entity s298 is
port (
G0: in std_logic; 
G1: in std_logic; 
G2: in std_logic; 
G117: out std_logic; 
G132: out std_logic; 
G66: out std_logic; 
G118: out std_logic; 
G133: out std_logic; 
G67: out std_logic 
);
end entity; 

architecture rtl of s298 is
begin
end architecture;
