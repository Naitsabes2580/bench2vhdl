--------------------------------------------------------------------------------
-- Testing signal G29 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G29;"));
signal_force("/s298_fc_tb/uut/G29", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G29", 0);
signal_force("/s298_fc_tb/uut/G29", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G29", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G10 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G10;"));
signal_force("/s298_fc_tb/uut/G10", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G10", 0);
signal_force("/s298_fc_tb/uut/G10", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G10", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G30 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G30;"));
signal_force("/s298_fc_tb/uut/G30", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G30", 0);
signal_force("/s298_fc_tb/uut/G30", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G30", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G11 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G11;"));
signal_force("/s298_fc_tb/uut/G11", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G11", 0);
signal_force("/s298_fc_tb/uut/G11", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G11", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G34 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G34;"));
signal_force("/s298_fc_tb/uut/G34", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G34", 0);
signal_force("/s298_fc_tb/uut/G34", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G34", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G12 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G12;"));
signal_force("/s298_fc_tb/uut/G12", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G12", 0);
signal_force("/s298_fc_tb/uut/G12", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G12", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G39 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G39;"));
signal_force("/s298_fc_tb/uut/G39", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G39", 0);
signal_force("/s298_fc_tb/uut/G39", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G39", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G13 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G13;"));
signal_force("/s298_fc_tb/uut/G13", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G13", 0);
signal_force("/s298_fc_tb/uut/G13", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G13", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G44 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G44;"));
signal_force("/s298_fc_tb/uut/G44", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G44", 0);
signal_force("/s298_fc_tb/uut/G44", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G44", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G14 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G14;"));
signal_force("/s298_fc_tb/uut/G14", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G14", 0);
signal_force("/s298_fc_tb/uut/G14", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G14", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G56 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G56;"));
signal_force("/s298_fc_tb/uut/G56", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G56", 0);
signal_force("/s298_fc_tb/uut/G56", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G56", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G15 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G15;"));
signal_force("/s298_fc_tb/uut/G15", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G15", 0);
signal_force("/s298_fc_tb/uut/G15", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G15", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G86 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G86;"));
signal_force("/s298_fc_tb/uut/G86", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G86", 0);
signal_force("/s298_fc_tb/uut/G86", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G86", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G16 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G16;"));
signal_force("/s298_fc_tb/uut/G16", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G16", 0);
signal_force("/s298_fc_tb/uut/G16", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G16", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G92 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G92;"));
signal_force("/s298_fc_tb/uut/G92", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G92", 0);
signal_force("/s298_fc_tb/uut/G92", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G92", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G17 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G17;"));
signal_force("/s298_fc_tb/uut/G17", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G17", 0);
signal_force("/s298_fc_tb/uut/G17", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G17", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G98 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G98;"));
signal_force("/s298_fc_tb/uut/G98", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G98", 0);
signal_force("/s298_fc_tb/uut/G98", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G98", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G18 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G18;"));
signal_force("/s298_fc_tb/uut/G18", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G18", 0);
signal_force("/s298_fc_tb/uut/G18", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G18", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G102 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G102;"));
signal_force("/s298_fc_tb/uut/G102", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G102", 0);
signal_force("/s298_fc_tb/uut/G102", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G102", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G19 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G19;"));
signal_force("/s298_fc_tb/uut/G19", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G19", 0);
signal_force("/s298_fc_tb/uut/G19", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G19", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G107 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G107;"));
signal_force("/s298_fc_tb/uut/G107", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G107", 0);
signal_force("/s298_fc_tb/uut/G107", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G107", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G20 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G20;"));
signal_force("/s298_fc_tb/uut/G20", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G20", 0);
signal_force("/s298_fc_tb/uut/G20", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G20", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G113 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G113;"));
signal_force("/s298_fc_tb/uut/G113", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G113", 0);
signal_force("/s298_fc_tb/uut/G113", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G113", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G21 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G21;"));
signal_force("/s298_fc_tb/uut/G21", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G21", 0);
signal_force("/s298_fc_tb/uut/G21", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G21", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G119 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G119;"));
signal_force("/s298_fc_tb/uut/G119", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G119", 0);
signal_force("/s298_fc_tb/uut/G119", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G119", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G22 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G22;"));
signal_force("/s298_fc_tb/uut/G22", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G22", 0);
signal_force("/s298_fc_tb/uut/G22", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G22", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G125 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G125;"));
signal_force("/s298_fc_tb/uut/G125", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G125", 0);
signal_force("/s298_fc_tb/uut/G125", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G125", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G23 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G23;"));
signal_force("/s298_fc_tb/uut/G23", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G23", 0);
signal_force("/s298_fc_tb/uut/G23", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G23", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G130 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G130;"));
signal_force("/s298_fc_tb/uut/G130", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G130", 0);
signal_force("/s298_fc_tb/uut/G130", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G130", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G28 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G28;"));
signal_force("/s298_fc_tb/uut/G28", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G28", 0);
signal_force("/s298_fc_tb/uut/G28", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G28", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G38 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G38;"));
signal_force("/s298_fc_tb/uut/G38", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G38", 0);
signal_force("/s298_fc_tb/uut/G38", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G38", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G40 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G40;"));
signal_force("/s298_fc_tb/uut/G40", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G40", 0);
signal_force("/s298_fc_tb/uut/G40", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G40", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G45 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G45;"));
signal_force("/s298_fc_tb/uut/G45", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G45", 0);
signal_force("/s298_fc_tb/uut/G45", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G45", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G46 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G46;"));
signal_force("/s298_fc_tb/uut/G46", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G46", 0);
signal_force("/s298_fc_tb/uut/G46", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G46", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G50 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G50;"));
signal_force("/s298_fc_tb/uut/G50", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G50", 0);
signal_force("/s298_fc_tb/uut/G50", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G50", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G51 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G51;"));
signal_force("/s298_fc_tb/uut/G51", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G51", 0);
signal_force("/s298_fc_tb/uut/G51", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G51", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G54 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G54;"));
signal_force("/s298_fc_tb/uut/G54", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G54", 0);
signal_force("/s298_fc_tb/uut/G54", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G54", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G55 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G55;"));
signal_force("/s298_fc_tb/uut/G55", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G55", 0);
signal_force("/s298_fc_tb/uut/G55", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G55", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G59 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G59;"));
signal_force("/s298_fc_tb/uut/G59", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G59", 0);
signal_force("/s298_fc_tb/uut/G59", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G59", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G60 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G60;"));
signal_force("/s298_fc_tb/uut/G60", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G60", 0);
signal_force("/s298_fc_tb/uut/G60", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G60", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G64 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G64;"));
signal_force("/s298_fc_tb/uut/G64", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G64", 0);
signal_force("/s298_fc_tb/uut/G64", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G64", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I155 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I155;"));
signal_force("/s298_fc_tb/uut/I155", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I155", 0);
signal_force("/s298_fc_tb/uut/I155", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I155", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I158 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I158;"));
signal_force("/s298_fc_tb/uut/I158", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I158", 0);
signal_force("/s298_fc_tb/uut/I158", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I158", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G76 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G76;"));
signal_force("/s298_fc_tb/uut/G76", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G76", 0);
signal_force("/s298_fc_tb/uut/G76", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G76", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G82 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G82;"));
signal_force("/s298_fc_tb/uut/G82", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G82", 0);
signal_force("/s298_fc_tb/uut/G82", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G82", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G87 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G87;"));
signal_force("/s298_fc_tb/uut/G87", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G87", 0);
signal_force("/s298_fc_tb/uut/G87", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G87", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G91 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G91;"));
signal_force("/s298_fc_tb/uut/G91", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G91", 0);
signal_force("/s298_fc_tb/uut/G91", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G91", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G93 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G93;"));
signal_force("/s298_fc_tb/uut/G93", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G93", 0);
signal_force("/s298_fc_tb/uut/G93", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G93", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G96 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G96;"));
signal_force("/s298_fc_tb/uut/G96", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G96", 0);
signal_force("/s298_fc_tb/uut/G96", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G96", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G99 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G99;"));
signal_force("/s298_fc_tb/uut/G99", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G99", 0);
signal_force("/s298_fc_tb/uut/G99", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G99", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G103 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G103;"));
signal_force("/s298_fc_tb/uut/G103", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G103", 0);
signal_force("/s298_fc_tb/uut/G103", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G103", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G112 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G112;"));
signal_force("/s298_fc_tb/uut/G112", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G112", 0);
signal_force("/s298_fc_tb/uut/G112", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G112", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G108 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G108;"));
signal_force("/s298_fc_tb/uut/G108", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G108", 0);
signal_force("/s298_fc_tb/uut/G108", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G108", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G114 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G114;"));
signal_force("/s298_fc_tb/uut/G114", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G114", 0);
signal_force("/s298_fc_tb/uut/G114", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G114", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I210 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I210;"));
signal_force("/s298_fc_tb/uut/I210", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I210", 0);
signal_force("/s298_fc_tb/uut/I210", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I210", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I213 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I213;"));
signal_force("/s298_fc_tb/uut/I213", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I213", 0);
signal_force("/s298_fc_tb/uut/I213", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I213", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G124 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G124;"));
signal_force("/s298_fc_tb/uut/G124", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G124", 0);
signal_force("/s298_fc_tb/uut/G124", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G124", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G120 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G120;"));
signal_force("/s298_fc_tb/uut/G120", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G120", 0);
signal_force("/s298_fc_tb/uut/G120", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G120", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G121 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G121;"));
signal_force("/s298_fc_tb/uut/G121", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G121", 0);
signal_force("/s298_fc_tb/uut/G121", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G121", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I221 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I221;"));
signal_force("/s298_fc_tb/uut/I221", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I221", 0);
signal_force("/s298_fc_tb/uut/I221", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I221", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G131 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G131;"));
signal_force("/s298_fc_tb/uut/G131", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G131", 0);
signal_force("/s298_fc_tb/uut/G131", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G131", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G126 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G126;"));
signal_force("/s298_fc_tb/uut/G126", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G126", 0);
signal_force("/s298_fc_tb/uut/G126", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G126", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G127 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G127;"));
signal_force("/s298_fc_tb/uut/G127", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G127", 0);
signal_force("/s298_fc_tb/uut/G127", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G127", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I229 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I229;"));
signal_force("/s298_fc_tb/uut/I229", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I229", 0);
signal_force("/s298_fc_tb/uut/I229", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I229", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I232 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I232;"));
signal_force("/s298_fc_tb/uut/I232", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I232", 0);
signal_force("/s298_fc_tb/uut/I232", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I232", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I235 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I235;"));
signal_force("/s298_fc_tb/uut/I235", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I235", 0);
signal_force("/s298_fc_tb/uut/I235", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I235", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I238 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I238;"));
signal_force("/s298_fc_tb/uut/I238", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I238", 0);
signal_force("/s298_fc_tb/uut/I238", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I238", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G26 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G26;"));
signal_force("/s298_fc_tb/uut/G26", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G26", 0);
signal_force("/s298_fc_tb/uut/G26", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G26", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G27 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G27;"));
signal_force("/s298_fc_tb/uut/G27", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G27", 0);
signal_force("/s298_fc_tb/uut/G27", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G27", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G31 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G31;"));
signal_force("/s298_fc_tb/uut/G31", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G31", 0);
signal_force("/s298_fc_tb/uut/G31", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G31", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G32 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G32;"));
signal_force("/s298_fc_tb/uut/G32", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G32", 0);
signal_force("/s298_fc_tb/uut/G32", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G32", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G33 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G33;"));
signal_force("/s298_fc_tb/uut/G33", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G33", 0);
signal_force("/s298_fc_tb/uut/G33", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G33", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G35 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G35;"));
signal_force("/s298_fc_tb/uut/G35", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G35", 0);
signal_force("/s298_fc_tb/uut/G35", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G35", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G36 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G36;"));
signal_force("/s298_fc_tb/uut/G36", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G36", 0);
signal_force("/s298_fc_tb/uut/G36", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G36", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G37 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G37;"));
signal_force("/s298_fc_tb/uut/G37", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G37", 0);
signal_force("/s298_fc_tb/uut/G37", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G37", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G42 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G42;"));
signal_force("/s298_fc_tb/uut/G42", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G42", 0);
signal_force("/s298_fc_tb/uut/G42", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G42", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G41 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G41;"));
signal_force("/s298_fc_tb/uut/G41", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G41", 0);
signal_force("/s298_fc_tb/uut/G41", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G41", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G48 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G48;"));
signal_force("/s298_fc_tb/uut/G48", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G48", 0);
signal_force("/s298_fc_tb/uut/G48", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G48", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G47 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G47;"));
signal_force("/s298_fc_tb/uut/G47", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G47", 0);
signal_force("/s298_fc_tb/uut/G47", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G47", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G49 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G49;"));
signal_force("/s298_fc_tb/uut/G49", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G49", 0);
signal_force("/s298_fc_tb/uut/G49", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G49", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G52 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G52;"));
signal_force("/s298_fc_tb/uut/G52", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G52", 0);
signal_force("/s298_fc_tb/uut/G52", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G52", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G57 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G57;"));
signal_force("/s298_fc_tb/uut/G57", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G57", 0);
signal_force("/s298_fc_tb/uut/G57", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G57", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G61 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G61;"));
signal_force("/s298_fc_tb/uut/G61", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G61", 0);
signal_force("/s298_fc_tb/uut/G61", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G61", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G58 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G58;"));
signal_force("/s298_fc_tb/uut/G58", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G58", 0);
signal_force("/s298_fc_tb/uut/G58", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G58", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G65 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G65;"));
signal_force("/s298_fc_tb/uut/G65", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G65", 0);
signal_force("/s298_fc_tb/uut/G65", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G65", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G62 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G62;"));
signal_force("/s298_fc_tb/uut/G62", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G62", 0);
signal_force("/s298_fc_tb/uut/G62", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G62", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G63 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G63;"));
signal_force("/s298_fc_tb/uut/G63", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G63", 0);
signal_force("/s298_fc_tb/uut/G63", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G63", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G74 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G74;"));
signal_force("/s298_fc_tb/uut/G74", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G74", 0);
signal_force("/s298_fc_tb/uut/G74", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G74", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G75 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G75;"));
signal_force("/s298_fc_tb/uut/G75", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G75", 0);
signal_force("/s298_fc_tb/uut/G75", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G75", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G88 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G88;"));
signal_force("/s298_fc_tb/uut/G88", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G88", 0);
signal_force("/s298_fc_tb/uut/G88", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G88", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G89 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G89;"));
signal_force("/s298_fc_tb/uut/G89", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G89", 0);
signal_force("/s298_fc_tb/uut/G89", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G89", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G90 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G90;"));
signal_force("/s298_fc_tb/uut/G90", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G90", 0);
signal_force("/s298_fc_tb/uut/G90", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G90", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G94 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G94;"));
signal_force("/s298_fc_tb/uut/G94", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G94", 0);
signal_force("/s298_fc_tb/uut/G94", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G94", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G95 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G95;"));
signal_force("/s298_fc_tb/uut/G95", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G95", 0);
signal_force("/s298_fc_tb/uut/G95", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G95", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G100 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G100;"));
signal_force("/s298_fc_tb/uut/G100", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G100", 0);
signal_force("/s298_fc_tb/uut/G100", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G100", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G105 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G105;"));
signal_force("/s298_fc_tb/uut/G105", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G105", 0);
signal_force("/s298_fc_tb/uut/G105", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G105", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G104 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G104;"));
signal_force("/s298_fc_tb/uut/G104", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G104", 0);
signal_force("/s298_fc_tb/uut/G104", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G104", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G110 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G110;"));
signal_force("/s298_fc_tb/uut/G110", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G110", 0);
signal_force("/s298_fc_tb/uut/G110", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G110", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G109 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G109;"));
signal_force("/s298_fc_tb/uut/G109", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G109", 0);
signal_force("/s298_fc_tb/uut/G109", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G109", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G111 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G111;"));
signal_force("/s298_fc_tb/uut/G111", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G111", 0);
signal_force("/s298_fc_tb/uut/G111", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G111", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G115 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G115;"));
signal_force("/s298_fc_tb/uut/G115", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G115", 0);
signal_force("/s298_fc_tb/uut/G115", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G115", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G122 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G122;"));
signal_force("/s298_fc_tb/uut/G122", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G122", 0);
signal_force("/s298_fc_tb/uut/G122", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G122", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G123 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G123;"));
signal_force("/s298_fc_tb/uut/G123", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G123", 0);
signal_force("/s298_fc_tb/uut/G123", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G123", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G128 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G128;"));
signal_force("/s298_fc_tb/uut/G128", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G128", 0);
signal_force("/s298_fc_tb/uut/G128", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G128", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G129 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G129;"));
signal_force("/s298_fc_tb/uut/G129", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G129", 0);
signal_force("/s298_fc_tb/uut/G129", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G129", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G24 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G24;"));
signal_force("/s298_fc_tb/uut/G24", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G24", 0);
signal_force("/s298_fc_tb/uut/G24", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G24", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G25 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G25;"));
signal_force("/s298_fc_tb/uut/G25", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G25", 0);
signal_force("/s298_fc_tb/uut/G25", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G25", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G68 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G68;"));
signal_force("/s298_fc_tb/uut/G68", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G68", 0);
signal_force("/s298_fc_tb/uut/G68", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G68", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G69 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G69;"));
signal_force("/s298_fc_tb/uut/G69", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G69", 0);
signal_force("/s298_fc_tb/uut/G69", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G69", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G70 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G70;"));
signal_force("/s298_fc_tb/uut/G70", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G70", 0);
signal_force("/s298_fc_tb/uut/G70", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G70", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G71 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G71;"));
signal_force("/s298_fc_tb/uut/G71", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G71", 0);
signal_force("/s298_fc_tb/uut/G71", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G71", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G72 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G72;"));
signal_force("/s298_fc_tb/uut/G72", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G72", 0);
signal_force("/s298_fc_tb/uut/G72", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G72", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G73 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G73;"));
signal_force("/s298_fc_tb/uut/G73", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G73", 0);
signal_force("/s298_fc_tb/uut/G73", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G73", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G77 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G77;"));
signal_force("/s298_fc_tb/uut/G77", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G77", 0);
signal_force("/s298_fc_tb/uut/G77", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G77", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G78 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G78;"));
signal_force("/s298_fc_tb/uut/G78", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G78", 0);
signal_force("/s298_fc_tb/uut/G78", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G78", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G79 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G79;"));
signal_force("/s298_fc_tb/uut/G79", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G79", 0);
signal_force("/s298_fc_tb/uut/G79", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G79", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G80 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G80;"));
signal_force("/s298_fc_tb/uut/G80", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G80", 0);
signal_force("/s298_fc_tb/uut/G80", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G80", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G81 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G81;"));
signal_force("/s298_fc_tb/uut/G81", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G81", 0);
signal_force("/s298_fc_tb/uut/G81", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G81", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G83 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G83;"));
signal_force("/s298_fc_tb/uut/G83", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G83", 0);
signal_force("/s298_fc_tb/uut/G83", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G83", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G84 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G84;"));
signal_force("/s298_fc_tb/uut/G84", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G84", 0);
signal_force("/s298_fc_tb/uut/G84", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G84", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G85 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G85;"));
signal_force("/s298_fc_tb/uut/G85", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G85", 0);
signal_force("/s298_fc_tb/uut/G85", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G85", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G43 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G43;"));
signal_force("/s298_fc_tb/uut/G43", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G43", 0);
signal_force("/s298_fc_tb/uut/G43", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G43", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G97 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G97;"));
signal_force("/s298_fc_tb/uut/G97", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G97", 0);
signal_force("/s298_fc_tb/uut/G97", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G97", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G101 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G101;"));
signal_force("/s298_fc_tb/uut/G101", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G101", 0);
signal_force("/s298_fc_tb/uut/G101", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G101", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G106 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G106;"));
signal_force("/s298_fc_tb/uut/G106", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G106", 0);
signal_force("/s298_fc_tb/uut/G106", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G106", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G116 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G116;"));
signal_force("/s298_fc_tb/uut/G116", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G116", 0);
signal_force("/s298_fc_tb/uut/G116", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G116", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G53 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G53;"));
signal_force("/s298_fc_tb/uut/G53", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G53", 0);
signal_force("/s298_fc_tb/uut/G53", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G53", 0);
writeline(out_file, s_a_line);
