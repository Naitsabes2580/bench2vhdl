--------------------------------------------------------------------------------
-- Testing signal G1 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G1;"));
signal_force("/s298_fc_tb/uut/G1", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G1", 0);
signal_force("/s298_fc_tb/uut/G1", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G1", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G2 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G2;"));
signal_force("/s298_fc_tb/uut/G2", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G2", 0);
signal_force("/s298_fc_tb/uut/G2", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G2", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G3 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G3;"));
signal_force("/s298_fc_tb/uut/G3", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G3", 0);
signal_force("/s298_fc_tb/uut/G3", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G3", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G4 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G4;"));
signal_force("/s298_fc_tb/uut/G4", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G4", 0);
signal_force("/s298_fc_tb/uut/G4", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G4", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G5 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G5;"));
signal_force("/s298_fc_tb/uut/G5", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G5", 0);
signal_force("/s298_fc_tb/uut/G5", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G5", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G6 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G6;"));
signal_force("/s298_fc_tb/uut/G6", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G6", 0);
signal_force("/s298_fc_tb/uut/G6", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G6", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G8 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G8;"));
signal_force("/s298_fc_tb/uut/G8", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G8", 0);
signal_force("/s298_fc_tb/uut/G8", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G8", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G9 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G9;"));
signal_force("/s298_fc_tb/uut/G9", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G9", 0);
signal_force("/s298_fc_tb/uut/G9", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G9", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G10 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G10;"));
signal_force("/s298_fc_tb/uut/G10", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G10", 0);
signal_force("/s298_fc_tb/uut/G10", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G10", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G11 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G11;"));
signal_force("/s298_fc_tb/uut/G11", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G11", 0);
signal_force("/s298_fc_tb/uut/G11", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G11", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G12 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G12;"));
signal_force("/s298_fc_tb/uut/G12", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G12", 0);
signal_force("/s298_fc_tb/uut/G12", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G12", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G13 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G13;"));
signal_force("/s298_fc_tb/uut/G13", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G13", 0);
signal_force("/s298_fc_tb/uut/G13", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G13", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G14 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G14;"));
signal_force("/s298_fc_tb/uut/G14", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G14", 0);
signal_force("/s298_fc_tb/uut/G14", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G14", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G15 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G15;"));
signal_force("/s298_fc_tb/uut/G15", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G15", 0);
signal_force("/s298_fc_tb/uut/G15", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G15", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G16 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G16;"));
signal_force("/s298_fc_tb/uut/G16", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G16", 0);
signal_force("/s298_fc_tb/uut/G16", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G16", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G17 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G17;"));
signal_force("/s298_fc_tb/uut/G17", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G17", 0);
signal_force("/s298_fc_tb/uut/G17", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G17", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G18 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G18;"));
signal_force("/s298_fc_tb/uut/G18", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G18", 0);
signal_force("/s298_fc_tb/uut/G18", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G18", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G19 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G19;"));
signal_force("/s298_fc_tb/uut/G19", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G19", 0);
signal_force("/s298_fc_tb/uut/G19", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G19", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G20 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G20;"));
signal_force("/s298_fc_tb/uut/G20", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G20", 0);
signal_force("/s298_fc_tb/uut/G20", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G20", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G21 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G21;"));
signal_force("/s298_fc_tb/uut/G21", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G21", 0);
signal_force("/s298_fc_tb/uut/G21", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G21", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G22 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G22;"));
signal_force("/s298_fc_tb/uut/G22", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G22", 0);
signal_force("/s298_fc_tb/uut/G22", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G22", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G23 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G23;"));
signal_force("/s298_fc_tb/uut/G23", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G23", 0);
signal_force("/s298_fc_tb/uut/G23", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G23", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G24 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G24;"));
signal_force("/s298_fc_tb/uut/G24", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G24", 0);
signal_force("/s298_fc_tb/uut/G24", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G24", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G25 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G25;"));
signal_force("/s298_fc_tb/uut/G25", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G25", 0);
signal_force("/s298_fc_tb/uut/G25", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G25", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G26 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G26;"));
signal_force("/s298_fc_tb/uut/G26", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G26", 0);
signal_force("/s298_fc_tb/uut/G26", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G26", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G27 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G27;"));
signal_force("/s298_fc_tb/uut/G27", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G27", 0);
signal_force("/s298_fc_tb/uut/G27", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G27", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G28 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G28;"));
signal_force("/s298_fc_tb/uut/G28", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G28", 0);
signal_force("/s298_fc_tb/uut/G28", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G28", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G29 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G29;"));
signal_force("/s298_fc_tb/uut/G29", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G29", 0);
signal_force("/s298_fc_tb/uut/G29", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G29", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G30 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G30;"));
signal_force("/s298_fc_tb/uut/G30", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G30", 0);
signal_force("/s298_fc_tb/uut/G30", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G30", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G31 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G31;"));
signal_force("/s298_fc_tb/uut/G31", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G31", 0);
signal_force("/s298_fc_tb/uut/G31", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G31", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G32 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G32;"));
signal_force("/s298_fc_tb/uut/G32", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G32", 0);
signal_force("/s298_fc_tb/uut/G32", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G32", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G33 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G33;"));
signal_force("/s298_fc_tb/uut/G33", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G33", 0);
signal_force("/s298_fc_tb/uut/G33", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G33", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G34 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G34;"));
signal_force("/s298_fc_tb/uut/G34", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G34", 0);
signal_force("/s298_fc_tb/uut/G34", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G34", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G35 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G35;"));
signal_force("/s298_fc_tb/uut/G35", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G35", 0);
signal_force("/s298_fc_tb/uut/G35", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G35", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G36 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G36;"));
signal_force("/s298_fc_tb/uut/G36", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G36", 0);
signal_force("/s298_fc_tb/uut/G36", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G36", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G103BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G103BF;"));
signal_force("/s298_fc_tb/uut/G103BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G103BF", 0);
signal_force("/s298_fc_tb/uut/G103BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G103BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G104BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G104BF;"));
signal_force("/s298_fc_tb/uut/G104BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G104BF", 0);
signal_force("/s298_fc_tb/uut/G104BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G104BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G105BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G105BF;"));
signal_force("/s298_fc_tb/uut/G105BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G105BF", 0);
signal_force("/s298_fc_tb/uut/G105BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G105BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G106BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G106BF;"));
signal_force("/s298_fc_tb/uut/G106BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G106BF", 0);
signal_force("/s298_fc_tb/uut/G106BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G106BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G107 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G107;"));
signal_force("/s298_fc_tb/uut/G107", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G107", 0);
signal_force("/s298_fc_tb/uut/G107", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G107", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G83 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G83;"));
signal_force("/s298_fc_tb/uut/G83", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G83", 0);
signal_force("/s298_fc_tb/uut/G83", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G83", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G84 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G84;"));
signal_force("/s298_fc_tb/uut/G84", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G84", 0);
signal_force("/s298_fc_tb/uut/G84", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G84", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G85 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G85;"));
signal_force("/s298_fc_tb/uut/G85", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G85", 0);
signal_force("/s298_fc_tb/uut/G85", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G85", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G86BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G86BF;"));
signal_force("/s298_fc_tb/uut/G86BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G86BF", 0);
signal_force("/s298_fc_tb/uut/G86BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G86BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G87BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G87BF;"));
signal_force("/s298_fc_tb/uut/G87BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G87BF", 0);
signal_force("/s298_fc_tb/uut/G87BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G87BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G88BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G88BF;"));
signal_force("/s298_fc_tb/uut/G88BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G88BF", 0);
signal_force("/s298_fc_tb/uut/G88BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G88BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G89BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G89BF;"));
signal_force("/s298_fc_tb/uut/G89BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G89BF", 0);
signal_force("/s298_fc_tb/uut/G89BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G89BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G90 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G90;"));
signal_force("/s298_fc_tb/uut/G90", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G90", 0);
signal_force("/s298_fc_tb/uut/G90", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G90", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G91 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G91;"));
signal_force("/s298_fc_tb/uut/G91", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G91", 0);
signal_force("/s298_fc_tb/uut/G91", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G91", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G92 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G92;"));
signal_force("/s298_fc_tb/uut/G92", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G92", 0);
signal_force("/s298_fc_tb/uut/G92", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G92", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G94 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G94;"));
signal_force("/s298_fc_tb/uut/G94", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G94", 0);
signal_force("/s298_fc_tb/uut/G94", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G94", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G95BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G95BF;"));
signal_force("/s298_fc_tb/uut/G95BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G95BF", 0);
signal_force("/s298_fc_tb/uut/G95BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G95BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G96BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G96BF;"));
signal_force("/s298_fc_tb/uut/G96BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G96BF", 0);
signal_force("/s298_fc_tb/uut/G96BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G96BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G97BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G97BF;"));
signal_force("/s298_fc_tb/uut/G97BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G97BF", 0);
signal_force("/s298_fc_tb/uut/G97BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G97BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G98BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G98BF;"));
signal_force("/s298_fc_tb/uut/G98BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G98BF", 0);
signal_force("/s298_fc_tb/uut/G98BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G98BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G99BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G99BF;"));
signal_force("/s298_fc_tb/uut/G99BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G99BF", 0);
signal_force("/s298_fc_tb/uut/G99BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G99BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G100BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G100BF;"));
signal_force("/s298_fc_tb/uut/G100BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G100BF", 0);
signal_force("/s298_fc_tb/uut/G100BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G100BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G101BF with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G101BF;"));
signal_force("/s298_fc_tb/uut/G101BF", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G101BF", 0);
signal_force("/s298_fc_tb/uut/G101BF", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G101BF", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G380 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G380;"));
signal_force("/s298_fc_tb/uut/G380", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G380", 0);
signal_force("/s298_fc_tb/uut/G380", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G380", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G64 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G64;"));
signal_force("/s298_fc_tb/uut/G64", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G64", 0);
signal_force("/s298_fc_tb/uut/G64", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G64", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G262 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G262;"));
signal_force("/s298_fc_tb/uut/G262", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G262", 0);
signal_force("/s298_fc_tb/uut/G262", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G262", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G65 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G65;"));
signal_force("/s298_fc_tb/uut/G65", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G65", 0);
signal_force("/s298_fc_tb/uut/G65", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G65", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G394 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G394;"));
signal_force("/s298_fc_tb/uut/G394", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G394", 0);
signal_force("/s298_fc_tb/uut/G394", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G394", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G66 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G66;"));
signal_force("/s298_fc_tb/uut/G66", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G66", 0);
signal_force("/s298_fc_tb/uut/G66", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G66", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G250 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G250;"));
signal_force("/s298_fc_tb/uut/G250", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G250", 0);
signal_force("/s298_fc_tb/uut/G250", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G250", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G67 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G67;"));
signal_force("/s298_fc_tb/uut/G67", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G67", 0);
signal_force("/s298_fc_tb/uut/G67", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G67", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G122 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G122;"));
signal_force("/s298_fc_tb/uut/G122", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G122", 0);
signal_force("/s298_fc_tb/uut/G122", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G122", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G68 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G68;"));
signal_force("/s298_fc_tb/uut/G68", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G68", 0);
signal_force("/s298_fc_tb/uut/G68", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G68", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G133 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G133;"));
signal_force("/s298_fc_tb/uut/G133", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G133", 0);
signal_force("/s298_fc_tb/uut/G133", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G133", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G69 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G69;"));
signal_force("/s298_fc_tb/uut/G69", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G69", 0);
signal_force("/s298_fc_tb/uut/G69", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G69", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G138 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G138;"));
signal_force("/s298_fc_tb/uut/G138", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G138", 0);
signal_force("/s298_fc_tb/uut/G138", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G138", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G70 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G70;"));
signal_force("/s298_fc_tb/uut/G70", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G70", 0);
signal_force("/s298_fc_tb/uut/G70", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G70", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G139 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G139;"));
signal_force("/s298_fc_tb/uut/G139", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G139", 0);
signal_force("/s298_fc_tb/uut/G139", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G139", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G71 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G71;"));
signal_force("/s298_fc_tb/uut/G71", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G71", 0);
signal_force("/s298_fc_tb/uut/G71", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G71", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G140 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G140;"));
signal_force("/s298_fc_tb/uut/G140", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G140", 0);
signal_force("/s298_fc_tb/uut/G140", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G140", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G72 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G72;"));
signal_force("/s298_fc_tb/uut/G72", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G72", 0);
signal_force("/s298_fc_tb/uut/G72", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G72", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G141 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G141;"));
signal_force("/s298_fc_tb/uut/G141", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G141", 0);
signal_force("/s298_fc_tb/uut/G141", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G141", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G73 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G73;"));
signal_force("/s298_fc_tb/uut/G73", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G73", 0);
signal_force("/s298_fc_tb/uut/G73", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G73", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G142 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G142;"));
signal_force("/s298_fc_tb/uut/G142", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G142", 0);
signal_force("/s298_fc_tb/uut/G142", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G142", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G74 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G74;"));
signal_force("/s298_fc_tb/uut/G74", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G74", 0);
signal_force("/s298_fc_tb/uut/G74", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G74", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G125 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G125;"));
signal_force("/s298_fc_tb/uut/G125", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G125", 0);
signal_force("/s298_fc_tb/uut/G125", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G125", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G75 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G75;"));
signal_force("/s298_fc_tb/uut/G75", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G75", 0);
signal_force("/s298_fc_tb/uut/G75", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G75", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G126 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G126;"));
signal_force("/s298_fc_tb/uut/G126", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G126", 0);
signal_force("/s298_fc_tb/uut/G126", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G126", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G76 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G76;"));
signal_force("/s298_fc_tb/uut/G76", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G76", 0);
signal_force("/s298_fc_tb/uut/G76", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G76", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G127 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G127;"));
signal_force("/s298_fc_tb/uut/G127", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G127", 0);
signal_force("/s298_fc_tb/uut/G127", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G127", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G77 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G77;"));
signal_force("/s298_fc_tb/uut/G77", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G77", 0);
signal_force("/s298_fc_tb/uut/G77", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G77", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G128 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G128;"));
signal_force("/s298_fc_tb/uut/G128", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G128", 0);
signal_force("/s298_fc_tb/uut/G128", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G128", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G78 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G78;"));
signal_force("/s298_fc_tb/uut/G78", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G78", 0);
signal_force("/s298_fc_tb/uut/G78", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G78", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G129 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G129;"));
signal_force("/s298_fc_tb/uut/G129", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G129", 0);
signal_force("/s298_fc_tb/uut/G129", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G129", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G79 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G79;"));
signal_force("/s298_fc_tb/uut/G79", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G79", 0);
signal_force("/s298_fc_tb/uut/G79", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G79", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G130 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G130;"));
signal_force("/s298_fc_tb/uut/G130", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G130", 0);
signal_force("/s298_fc_tb/uut/G130", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G130", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G80 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G80;"));
signal_force("/s298_fc_tb/uut/G80", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G80", 0);
signal_force("/s298_fc_tb/uut/G80", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G80", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G131 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G131;"));
signal_force("/s298_fc_tb/uut/G131", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G131", 0);
signal_force("/s298_fc_tb/uut/G131", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G131", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G81 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G81;"));
signal_force("/s298_fc_tb/uut/G81", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G81", 0);
signal_force("/s298_fc_tb/uut/G81", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G81", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G132 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G132;"));
signal_force("/s298_fc_tb/uut/G132", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G132", 0);
signal_force("/s298_fc_tb/uut/G132", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G132", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G82 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G82;"));
signal_force("/s298_fc_tb/uut/G82", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G82", 0);
signal_force("/s298_fc_tb/uut/G82", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G82", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I633 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I633;"));
signal_force("/s298_fc_tb/uut/I633", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I633", 0);
signal_force("/s298_fc_tb/uut/I633", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I633", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G366 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G366;"));
signal_force("/s298_fc_tb/uut/G366", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G366", 0);
signal_force("/s298_fc_tb/uut/G366", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G366", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G379 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G379;"));
signal_force("/s298_fc_tb/uut/G379", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G379", 0);
signal_force("/s298_fc_tb/uut/G379", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G379", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I643 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I643;"));
signal_force("/s298_fc_tb/uut/I643", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I643", 0);
signal_force("/s298_fc_tb/uut/I643", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I643", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I646 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I646;"));
signal_force("/s298_fc_tb/uut/I646", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I646", 0);
signal_force("/s298_fc_tb/uut/I646", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I646", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I649 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I649;"));
signal_force("/s298_fc_tb/uut/I649", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I649", 0);
signal_force("/s298_fc_tb/uut/I649", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I649", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I652 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I652;"));
signal_force("/s298_fc_tb/uut/I652", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I652", 0);
signal_force("/s298_fc_tb/uut/I652", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I652", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I655 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I655;"));
signal_force("/s298_fc_tb/uut/I655", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I655", 0);
signal_force("/s298_fc_tb/uut/I655", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I655", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I660 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I660;"));
signal_force("/s298_fc_tb/uut/I660", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I660", 0);
signal_force("/s298_fc_tb/uut/I660", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I660", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I680 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I680;"));
signal_force("/s298_fc_tb/uut/I680", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I680", 0);
signal_force("/s298_fc_tb/uut/I680", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I680", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I684 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I684;"));
signal_force("/s298_fc_tb/uut/I684", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I684", 0);
signal_force("/s298_fc_tb/uut/I684", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I684", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I687 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I687;"));
signal_force("/s298_fc_tb/uut/I687", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I687", 0);
signal_force("/s298_fc_tb/uut/I687", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I687", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I165 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I165;"));
signal_force("/s298_fc_tb/uut/I165", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I165", 0);
signal_force("/s298_fc_tb/uut/I165", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I165", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G29 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G29;"));
signal_force("/s298_fc_tb/uut/G29", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G29", 0);
signal_force("/s298_fc_tb/uut/G29", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G29", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II178 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II178;"));
signal_force("/s298_fc_tb/uut/II178", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II178", 0);
signal_force("/s298_fc_tb/uut/II178", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II178", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I169 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I169;"));
signal_force("/s298_fc_tb/uut/I169", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I169", 0);
signal_force("/s298_fc_tb/uut/I169", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I169", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G113 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G113;"));
signal_force("/s298_fc_tb/uut/G113", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G113", 0);
signal_force("/s298_fc_tb/uut/G113", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G113", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I172 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I172;"));
signal_force("/s298_fc_tb/uut/I172", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I172", 0);
signal_force("/s298_fc_tb/uut/I172", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I172", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G115 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G115;"));
signal_force("/s298_fc_tb/uut/G115", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G115", 0);
signal_force("/s298_fc_tb/uut/G115", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G115", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I175 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I175;"));
signal_force("/s298_fc_tb/uut/I175", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I175", 0);
signal_force("/s298_fc_tb/uut/I175", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I175", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G117 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G117;"));
signal_force("/s298_fc_tb/uut/G117", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G117", 0);
signal_force("/s298_fc_tb/uut/G117", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G117", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I178 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I178;"));
signal_force("/s298_fc_tb/uut/I178", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I178", 0);
signal_force("/s298_fc_tb/uut/I178", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I178", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G219 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G219;"));
signal_force("/s298_fc_tb/uut/G219", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G219", 0);
signal_force("/s298_fc_tb/uut/G219", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G219", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I181 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I181;"));
signal_force("/s298_fc_tb/uut/I181", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I181", 0);
signal_force("/s298_fc_tb/uut/I181", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I181", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G119 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G119;"));
signal_force("/s298_fc_tb/uut/G119", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G119", 0);
signal_force("/s298_fc_tb/uut/G119", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G119", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I184 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I184;"));
signal_force("/s298_fc_tb/uut/I184", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I184", 0);
signal_force("/s298_fc_tb/uut/I184", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I184", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G221 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G221;"));
signal_force("/s298_fc_tb/uut/G221", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G221", 0);
signal_force("/s298_fc_tb/uut/G221", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G221", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I187 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I187;"));
signal_force("/s298_fc_tb/uut/I187", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I187", 0);
signal_force("/s298_fc_tb/uut/I187", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I187", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G121 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G121;"));
signal_force("/s298_fc_tb/uut/G121", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G121", 0);
signal_force("/s298_fc_tb/uut/G121", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G121", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I190 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I190;"));
signal_force("/s298_fc_tb/uut/I190", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I190", 0);
signal_force("/s298_fc_tb/uut/I190", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I190", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G223 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G223;"));
signal_force("/s298_fc_tb/uut/G223", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G223", 0);
signal_force("/s298_fc_tb/uut/G223", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G223", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I193 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I193;"));
signal_force("/s298_fc_tb/uut/I193", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I193", 0);
signal_force("/s298_fc_tb/uut/I193", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I193", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G209 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G209;"));
signal_force("/s298_fc_tb/uut/G209", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G209", 0);
signal_force("/s298_fc_tb/uut/G209", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G209", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I196 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I196;"));
signal_force("/s298_fc_tb/uut/I196", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I196", 0);
signal_force("/s298_fc_tb/uut/I196", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I196", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G109 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G109;"));
signal_force("/s298_fc_tb/uut/G109", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G109", 0);
signal_force("/s298_fc_tb/uut/G109", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G109", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I199 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I199;"));
signal_force("/s298_fc_tb/uut/I199", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I199", 0);
signal_force("/s298_fc_tb/uut/I199", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I199", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G211 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G211;"));
signal_force("/s298_fc_tb/uut/G211", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G211", 0);
signal_force("/s298_fc_tb/uut/G211", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G211", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I202 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I202;"));
signal_force("/s298_fc_tb/uut/I202", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I202", 0);
signal_force("/s298_fc_tb/uut/I202", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I202", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G111 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G111;"));
signal_force("/s298_fc_tb/uut/G111", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G111", 0);
signal_force("/s298_fc_tb/uut/G111", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G111", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I205 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I205;"));
signal_force("/s298_fc_tb/uut/I205", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I205", 0);
signal_force("/s298_fc_tb/uut/I205", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I205", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G213 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G213;"));
signal_force("/s298_fc_tb/uut/G213", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G213", 0);
signal_force("/s298_fc_tb/uut/G213", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G213", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I208 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I208;"));
signal_force("/s298_fc_tb/uut/I208", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I208", 0);
signal_force("/s298_fc_tb/uut/I208", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I208", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G215 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G215;"));
signal_force("/s298_fc_tb/uut/G215", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G215", 0);
signal_force("/s298_fc_tb/uut/G215", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G215", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I211 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I211;"));
signal_force("/s298_fc_tb/uut/I211", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I211", 0);
signal_force("/s298_fc_tb/uut/I211", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I211", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G217 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G217;"));
signal_force("/s298_fc_tb/uut/G217", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G217", 0);
signal_force("/s298_fc_tb/uut/G217", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G217", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G352 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G352;"));
signal_force("/s298_fc_tb/uut/G352", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G352", 0);
signal_force("/s298_fc_tb/uut/G352", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G352", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G360 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G360;"));
signal_force("/s298_fc_tb/uut/G360", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G360", 0);
signal_force("/s298_fc_tb/uut/G360", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G360", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G361 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G361;"));
signal_force("/s298_fc_tb/uut/G361", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G361", 0);
signal_force("/s298_fc_tb/uut/G361", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G361", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G362 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G362;"));
signal_force("/s298_fc_tb/uut/G362", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G362", 0);
signal_force("/s298_fc_tb/uut/G362", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G362", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G363 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G363;"));
signal_force("/s298_fc_tb/uut/G363", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G363", 0);
signal_force("/s298_fc_tb/uut/G363", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G363", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G364 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G364;"));
signal_force("/s298_fc_tb/uut/G364", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G364", 0);
signal_force("/s298_fc_tb/uut/G364", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G364", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G367 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G367;"));
signal_force("/s298_fc_tb/uut/G367", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G367", 0);
signal_force("/s298_fc_tb/uut/G367", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G367", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G386 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G386;"));
signal_force("/s298_fc_tb/uut/G386", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G386", 0);
signal_force("/s298_fc_tb/uut/G386", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G386", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G388 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G388;"));
signal_force("/s298_fc_tb/uut/G388", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G388", 0);
signal_force("/s298_fc_tb/uut/G388", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G388", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G389 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G389;"));
signal_force("/s298_fc_tb/uut/G389", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G389", 0);
signal_force("/s298_fc_tb/uut/G389", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G389", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G110 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G110;"));
signal_force("/s298_fc_tb/uut/G110", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G110", 0);
signal_force("/s298_fc_tb/uut/G110", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G110", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G114 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G114;"));
signal_force("/s298_fc_tb/uut/G114", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G114", 0);
signal_force("/s298_fc_tb/uut/G114", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G114", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G118 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G118;"));
signal_force("/s298_fc_tb/uut/G118", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G118", 0);
signal_force("/s298_fc_tb/uut/G118", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G118", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G216 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G216;"));
signal_force("/s298_fc_tb/uut/G216", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G216", 0);
signal_force("/s298_fc_tb/uut/G216", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G216", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G218 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G218;"));
signal_force("/s298_fc_tb/uut/G218", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G218", 0);
signal_force("/s298_fc_tb/uut/G218", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G218", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G220 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G220;"));
signal_force("/s298_fc_tb/uut/G220", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G220", 0);
signal_force("/s298_fc_tb/uut/G220", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G220", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G222 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G222;"));
signal_force("/s298_fc_tb/uut/G222", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G222", 0);
signal_force("/s298_fc_tb/uut/G222", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G222", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G365 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G365;"));
signal_force("/s298_fc_tb/uut/G365", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G365", 0);
signal_force("/s298_fc_tb/uut/G365", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G365", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G368 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G368;"));
signal_force("/s298_fc_tb/uut/G368", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G368", 0);
signal_force("/s298_fc_tb/uut/G368", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G368", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G387 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G387;"));
signal_force("/s298_fc_tb/uut/G387", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G387", 0);
signal_force("/s298_fc_tb/uut/G387", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G387", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G225 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G225;"));
signal_force("/s298_fc_tb/uut/G225", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G225", 0);
signal_force("/s298_fc_tb/uut/G225", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G225", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G390 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G390;"));
signal_force("/s298_fc_tb/uut/G390", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G390", 0);
signal_force("/s298_fc_tb/uut/G390", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G390", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G289 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G289;"));
signal_force("/s298_fc_tb/uut/G289", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G289", 0);
signal_force("/s298_fc_tb/uut/G289", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G289", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I356 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I356;"));
signal_force("/s298_fc_tb/uut/I356", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I356", 0);
signal_force("/s298_fc_tb/uut/I356", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I356", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G324 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G324;"));
signal_force("/s298_fc_tb/uut/G324", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G324", 0);
signal_force("/s298_fc_tb/uut/G324", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G324", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I254 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I254;"));
signal_force("/s298_fc_tb/uut/I254", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I254", 0);
signal_force("/s298_fc_tb/uut/I254", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I254", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G166 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G166;"));
signal_force("/s298_fc_tb/uut/G166", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G166", 0);
signal_force("/s298_fc_tb/uut/G166", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G166", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I257 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I257;"));
signal_force("/s298_fc_tb/uut/I257", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I257", 0);
signal_force("/s298_fc_tb/uut/I257", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I257", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G325 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G325;"));
signal_force("/s298_fc_tb/uut/G325", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G325", 0);
signal_force("/s298_fc_tb/uut/G325", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G325", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G338 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G338;"));
signal_force("/s298_fc_tb/uut/G338", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G338", 0);
signal_force("/s298_fc_tb/uut/G338", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G338", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I260 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I260;"));
signal_force("/s298_fc_tb/uut/I260", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I260", 0);
signal_force("/s298_fc_tb/uut/I260", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I260", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G194 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G194;"));
signal_force("/s298_fc_tb/uut/G194", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G194", 0);
signal_force("/s298_fc_tb/uut/G194", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G194", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I263 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I263;"));
signal_force("/s298_fc_tb/uut/I263", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I263", 0);
signal_force("/s298_fc_tb/uut/I263", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I263", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G339 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G339;"));
signal_force("/s298_fc_tb/uut/G339", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G339", 0);
signal_force("/s298_fc_tb/uut/G339", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G339", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G344 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G344;"));
signal_force("/s298_fc_tb/uut/G344", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G344", 0);
signal_force("/s298_fc_tb/uut/G344", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G344", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I266 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I266;"));
signal_force("/s298_fc_tb/uut/I266", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I266", 0);
signal_force("/s298_fc_tb/uut/I266", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I266", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G202 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G202;"));
signal_force("/s298_fc_tb/uut/G202", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G202", 0);
signal_force("/s298_fc_tb/uut/G202", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G202", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I269 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I269;"));
signal_force("/s298_fc_tb/uut/I269", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I269", 0);
signal_force("/s298_fc_tb/uut/I269", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I269", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G345 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G345;"));
signal_force("/s298_fc_tb/uut/G345", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G345", 0);
signal_force("/s298_fc_tb/uut/G345", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G345", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G312 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G312;"));
signal_force("/s298_fc_tb/uut/G312", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G312", 0);
signal_force("/s298_fc_tb/uut/G312", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G312", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I272 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I272;"));
signal_force("/s298_fc_tb/uut/I272", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I272", 0);
signal_force("/s298_fc_tb/uut/I272", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I272", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G313 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G313;"));
signal_force("/s298_fc_tb/uut/G313", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G313", 0);
signal_force("/s298_fc_tb/uut/G313", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G313", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G315 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G315;"));
signal_force("/s298_fc_tb/uut/G315", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G315", 0);
signal_force("/s298_fc_tb/uut/G315", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G315", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I275 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I275;"));
signal_force("/s298_fc_tb/uut/I275", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I275", 0);
signal_force("/s298_fc_tb/uut/I275", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I275", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G316 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G316;"));
signal_force("/s298_fc_tb/uut/G316", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G316", 0);
signal_force("/s298_fc_tb/uut/G316", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G316", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G318 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G318;"));
signal_force("/s298_fc_tb/uut/G318", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G318", 0);
signal_force("/s298_fc_tb/uut/G318", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G318", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I278 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I278;"));
signal_force("/s298_fc_tb/uut/I278", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I278", 0);
signal_force("/s298_fc_tb/uut/I278", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I278", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G319 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G319;"));
signal_force("/s298_fc_tb/uut/G319", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G319", 0);
signal_force("/s298_fc_tb/uut/G319", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G319", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G321 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G321;"));
signal_force("/s298_fc_tb/uut/G321", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G321", 0);
signal_force("/s298_fc_tb/uut/G321", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G321", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I281 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I281;"));
signal_force("/s298_fc_tb/uut/I281", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I281", 0);
signal_force("/s298_fc_tb/uut/I281", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I281", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G322 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G322;"));
signal_force("/s298_fc_tb/uut/G322", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G322", 0);
signal_force("/s298_fc_tb/uut/G322", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G322", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G143 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G143;"));
signal_force("/s298_fc_tb/uut/G143", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G143", 0);
signal_force("/s298_fc_tb/uut/G143", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G143", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I287 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I287;"));
signal_force("/s298_fc_tb/uut/I287", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I287", 0);
signal_force("/s298_fc_tb/uut/I287", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I287", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G381 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G381;"));
signal_force("/s298_fc_tb/uut/G381", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G381", 0);
signal_force("/s298_fc_tb/uut/G381", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G381", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I291 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I291;"));
signal_force("/s298_fc_tb/uut/I291", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I291", 0);
signal_force("/s298_fc_tb/uut/I291", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I291", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G375 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G375;"));
signal_force("/s298_fc_tb/uut/G375", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G375", 0);
signal_force("/s298_fc_tb/uut/G375", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G375", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I295 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I295;"));
signal_force("/s298_fc_tb/uut/I295", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I295", 0);
signal_force("/s298_fc_tb/uut/I295", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I295", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G371 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G371;"));
signal_force("/s298_fc_tb/uut/G371", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G371", 0);
signal_force("/s298_fc_tb/uut/G371", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G371", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I303 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I303;"));
signal_force("/s298_fc_tb/uut/I303", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I303", 0);
signal_force("/s298_fc_tb/uut/I303", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I303", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G350 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G350;"));
signal_force("/s298_fc_tb/uut/G350", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G350", 0);
signal_force("/s298_fc_tb/uut/G350", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G350", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G281 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G281;"));
signal_force("/s298_fc_tb/uut/G281", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G281", 0);
signal_force("/s298_fc_tb/uut/G281", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G281", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I299 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I299;"));
signal_force("/s298_fc_tb/uut/I299", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I299", 0);
signal_force("/s298_fc_tb/uut/I299", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I299", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G283 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G283;"));
signal_force("/s298_fc_tb/uut/G283", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G283", 0);
signal_force("/s298_fc_tb/uut/G283", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G283", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I313 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I313;"));
signal_force("/s298_fc_tb/uut/I313", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I313", 0);
signal_force("/s298_fc_tb/uut/I313", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I313", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G382 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G382;"));
signal_force("/s298_fc_tb/uut/G382", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G382", 0);
signal_force("/s298_fc_tb/uut/G382", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G382", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G100 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G100;"));
signal_force("/s298_fc_tb/uut/G100", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G100", 0);
signal_force("/s298_fc_tb/uut/G100", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G100", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G376 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G376;"));
signal_force("/s298_fc_tb/uut/G376", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G376", 0);
signal_force("/s298_fc_tb/uut/G376", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G376", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G98 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G98;"));
signal_force("/s298_fc_tb/uut/G98", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G98", 0);
signal_force("/s298_fc_tb/uut/G98", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G98", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G372 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G372;"));
signal_force("/s298_fc_tb/uut/G372", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G372", 0);
signal_force("/s298_fc_tb/uut/G372", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G372", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G96 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G96;"));
signal_force("/s298_fc_tb/uut/G96", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G96", 0);
signal_force("/s298_fc_tb/uut/G96", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G96", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I301 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I301;"));
signal_force("/s298_fc_tb/uut/I301", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I301", 0);
signal_force("/s298_fc_tb/uut/I301", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I301", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I315 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I315;"));
signal_force("/s298_fc_tb/uut/I315", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I315", 0);
signal_force("/s298_fc_tb/uut/I315", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I315", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G135 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G135;"));
signal_force("/s298_fc_tb/uut/G135", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G135", 0);
signal_force("/s298_fc_tb/uut/G135", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G135", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I321 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I321;"));
signal_force("/s298_fc_tb/uut/I321", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I321", 0);
signal_force("/s298_fc_tb/uut/I321", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I321", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G329 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G329;"));
signal_force("/s298_fc_tb/uut/G329", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G329", 0);
signal_force("/s298_fc_tb/uut/G329", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G329", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G137 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G137;"));
signal_force("/s298_fc_tb/uut/G137", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G137", 0);
signal_force("/s298_fc_tb/uut/G137", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G137", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I324 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I324;"));
signal_force("/s298_fc_tb/uut/I324", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I324", 0);
signal_force("/s298_fc_tb/uut/I324", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I324", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G333 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G333;"));
signal_force("/s298_fc_tb/uut/G333", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G333", 0);
signal_force("/s298_fc_tb/uut/G333", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G333", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G87 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G87;"));
signal_force("/s298_fc_tb/uut/G87", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G87", 0);
signal_force("/s298_fc_tb/uut/G87", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G87", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I406 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I406;"));
signal_force("/s298_fc_tb/uut/I406", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I406", 0);
signal_force("/s298_fc_tb/uut/I406", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I406", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G89 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G89;"));
signal_force("/s298_fc_tb/uut/G89", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G89", 0);
signal_force("/s298_fc_tb/uut/G89", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G89", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I422 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I422;"));
signal_force("/s298_fc_tb/uut/I422", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I422", 0);
signal_force("/s298_fc_tb/uut/I422", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I422", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G173 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G173;"));
signal_force("/s298_fc_tb/uut/G173", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G173", 0);
signal_force("/s298_fc_tb/uut/G173", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G173", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G183 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G183;"));
signal_force("/s298_fc_tb/uut/G183", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G183", 0);
signal_force("/s298_fc_tb/uut/G183", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G183", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I335 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I335;"));
signal_force("/s298_fc_tb/uut/I335", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I335", 0);
signal_force("/s298_fc_tb/uut/I335", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I335", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G174 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G174;"));
signal_force("/s298_fc_tb/uut/G174", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G174", 0);
signal_force("/s298_fc_tb/uut/G174", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G174", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I338 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I338;"));
signal_force("/s298_fc_tb/uut/I338", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I338", 0);
signal_force("/s298_fc_tb/uut/I338", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I338", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G184 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G184;"));
signal_force("/s298_fc_tb/uut/G184", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G184", 0);
signal_force("/s298_fc_tb/uut/G184", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G184", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I341 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I341;"));
signal_force("/s298_fc_tb/uut/I341", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I341", 0);
signal_force("/s298_fc_tb/uut/I341", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I341", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G355 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G355;"));
signal_force("/s298_fc_tb/uut/G355", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G355", 0);
signal_force("/s298_fc_tb/uut/G355", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G355", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G359 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G359;"));
signal_force("/s298_fc_tb/uut/G359", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G359", 0);
signal_force("/s298_fc_tb/uut/G359", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G359", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G356 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G356;"));
signal_force("/s298_fc_tb/uut/G356", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G356", 0);
signal_force("/s298_fc_tb/uut/G356", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G356", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G108 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G108;"));
signal_force("/s298_fc_tb/uut/G108", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G108", 0);
signal_force("/s298_fc_tb/uut/G108", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G108", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G116 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G116;"));
signal_force("/s298_fc_tb/uut/G116", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G116", 0);
signal_force("/s298_fc_tb/uut/G116", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G116", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G293 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G293;"));
signal_force("/s298_fc_tb/uut/G293", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G293", 0);
signal_force("/s298_fc_tb/uut/G293", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G293", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I354 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I354;"));
signal_force("/s298_fc_tb/uut/I354", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I354", 0);
signal_force("/s298_fc_tb/uut/I354", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I354", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G146 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G146;"));
signal_force("/s298_fc_tb/uut/G146", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G146", 0);
signal_force("/s298_fc_tb/uut/G146", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G146", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I357 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I357;"));
signal_force("/s298_fc_tb/uut/I357", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I357", 0);
signal_force("/s298_fc_tb/uut/I357", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I357", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G294 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G294;"));
signal_force("/s298_fc_tb/uut/G294", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G294", 0);
signal_force("/s298_fc_tb/uut/G294", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G294", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G309 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G309;"));
signal_force("/s298_fc_tb/uut/G309", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G309", 0);
signal_force("/s298_fc_tb/uut/G309", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G309", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I360 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I360;"));
signal_force("/s298_fc_tb/uut/I360", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I360", 0);
signal_force("/s298_fc_tb/uut/I360", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I360", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G162 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G162;"));
signal_force("/s298_fc_tb/uut/G162", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G162", 0);
signal_force("/s298_fc_tb/uut/G162", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G162", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I363 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I363;"));
signal_force("/s298_fc_tb/uut/I363", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I363", 0);
signal_force("/s298_fc_tb/uut/I363", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I363", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G310 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G310;"));
signal_force("/s298_fc_tb/uut/G310", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G310", 0);
signal_force("/s298_fc_tb/uut/G310", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G310", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G341 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G341;"));
signal_force("/s298_fc_tb/uut/G341", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G341", 0);
signal_force("/s298_fc_tb/uut/G341", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G341", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I366 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I366;"));
signal_force("/s298_fc_tb/uut/I366", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I366", 0);
signal_force("/s298_fc_tb/uut/I366", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I366", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G198 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G198;"));
signal_force("/s298_fc_tb/uut/G198", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G198", 0);
signal_force("/s298_fc_tb/uut/G198", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G198", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I369 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I369;"));
signal_force("/s298_fc_tb/uut/I369", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I369", 0);
signal_force("/s298_fc_tb/uut/I369", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I369", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G342 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G342;"));
signal_force("/s298_fc_tb/uut/G342", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G342", 0);
signal_force("/s298_fc_tb/uut/G342", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G342", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G303 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G303;"));
signal_force("/s298_fc_tb/uut/G303", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G303", 0);
signal_force("/s298_fc_tb/uut/G303", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G303", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I372 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I372;"));
signal_force("/s298_fc_tb/uut/I372", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I372", 0);
signal_force("/s298_fc_tb/uut/I372", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I372", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G154 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G154;"));
signal_force("/s298_fc_tb/uut/G154", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G154", 0);
signal_force("/s298_fc_tb/uut/G154", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G154", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I375 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I375;"));
signal_force("/s298_fc_tb/uut/I375", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I375", 0);
signal_force("/s298_fc_tb/uut/I375", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I375", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G304 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G304;"));
signal_force("/s298_fc_tb/uut/G304", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G304", 0);
signal_force("/s298_fc_tb/uut/G304", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G304", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I378 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I378;"));
signal_force("/s298_fc_tb/uut/I378", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I378", 0);
signal_force("/s298_fc_tb/uut/I378", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I378", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G383 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G383;"));
signal_force("/s298_fc_tb/uut/G383", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G383", 0);
signal_force("/s298_fc_tb/uut/G383", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G383", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I382 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I382;"));
signal_force("/s298_fc_tb/uut/I382", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I382", 0);
signal_force("/s298_fc_tb/uut/I382", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I382", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G396 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G396;"));
signal_force("/s298_fc_tb/uut/G396", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G396", 0);
signal_force("/s298_fc_tb/uut/G396", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G396", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I386 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I386;"));
signal_force("/s298_fc_tb/uut/I386", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I386", 0);
signal_force("/s298_fc_tb/uut/I386", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I386", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G373 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G373;"));
signal_force("/s298_fc_tb/uut/G373", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G373", 0);
signal_force("/s298_fc_tb/uut/G373", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G373", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I390 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I390;"));
signal_force("/s298_fc_tb/uut/I390", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I390", 0);
signal_force("/s298_fc_tb/uut/I390", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I390", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G392 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G392;"));
signal_force("/s298_fc_tb/uut/G392", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G392", 0);
signal_force("/s298_fc_tb/uut/G392", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G392", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G384 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G384;"));
signal_force("/s298_fc_tb/uut/G384", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G384", 0);
signal_force("/s298_fc_tb/uut/G384", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G384", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G101 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G101;"));
signal_force("/s298_fc_tb/uut/G101", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G101", 0);
signal_force("/s298_fc_tb/uut/G101", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G101", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G397 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G397;"));
signal_force("/s298_fc_tb/uut/G397", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G397", 0);
signal_force("/s298_fc_tb/uut/G397", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G397", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G106 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G106;"));
signal_force("/s298_fc_tb/uut/G106", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G106", 0);
signal_force("/s298_fc_tb/uut/G106", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G106", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G374 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G374;"));
signal_force("/s298_fc_tb/uut/G374", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G374", 0);
signal_force("/s298_fc_tb/uut/G374", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G374", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G97 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G97;"));
signal_force("/s298_fc_tb/uut/G97", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G97", 0);
signal_force("/s298_fc_tb/uut/G97", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G97", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G393 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G393;"));
signal_force("/s298_fc_tb/uut/G393", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G393", 0);
signal_force("/s298_fc_tb/uut/G393", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G393", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G104 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G104;"));
signal_force("/s298_fc_tb/uut/G104", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G104", 0);
signal_force("/s298_fc_tb/uut/G104", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G104", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II476 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II476;"));
signal_force("/s298_fc_tb/uut/II476", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II476", 0);
signal_force("/s298_fc_tb/uut/II476", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II476", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G278 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G278;"));
signal_force("/s298_fc_tb/uut/G278", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G278", 0);
signal_force("/s298_fc_tb/uut/G278", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G278", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I279 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I279;"));
signal_force("/s298_fc_tb/uut/I279", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I279", 0);
signal_force("/s298_fc_tb/uut/I279", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I279", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G224 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G224;"));
signal_force("/s298_fc_tb/uut/G224", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G224", 0);
signal_force("/s298_fc_tb/uut/G224", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G224", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G282 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G282;"));
signal_force("/s298_fc_tb/uut/G282", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G282", 0);
signal_force("/s298_fc_tb/uut/G282", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G282", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I306 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I306;"));
signal_force("/s298_fc_tb/uut/I306", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I306", 0);
signal_force("/s298_fc_tb/uut/I306", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I306", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G286 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G286;"));
signal_force("/s298_fc_tb/uut/G286", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G286", 0);
signal_force("/s298_fc_tb/uut/G286", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G286", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I334 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I334;"));
signal_force("/s298_fc_tb/uut/I334", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I334", 0);
signal_force("/s298_fc_tb/uut/I334", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I334", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G285 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G285;"));
signal_force("/s298_fc_tb/uut/G285", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G285", 0);
signal_force("/s298_fc_tb/uut/G285", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G285", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I327 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I327;"));
signal_force("/s298_fc_tb/uut/I327", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I327", 0);
signal_force("/s298_fc_tb/uut/I327", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I327", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G268 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G268;"));
signal_force("/s298_fc_tb/uut/G268", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G268", 0);
signal_force("/s298_fc_tb/uut/G268", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G268", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II208 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II208;"));
signal_force("/s298_fc_tb/uut/II208", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II208", 0);
signal_force("/s298_fc_tb/uut/II208", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II208", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I308 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I308;"));
signal_force("/s298_fc_tb/uut/I308", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I308", 0);
signal_force("/s298_fc_tb/uut/I308", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I308", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I336 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I336;"));
signal_force("/s298_fc_tb/uut/I336", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I336", 0);
signal_force("/s298_fc_tb/uut/I336", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I336", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I329 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I329;"));
signal_force("/s298_fc_tb/uut/I329", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I329", 0);
signal_force("/s298_fc_tb/uut/I329", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I329", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I210 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I210;"));
signal_force("/s298_fc_tb/uut/I210", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I210", 0);
signal_force("/s298_fc_tb/uut/I210", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I210", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G136 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G136;"));
signal_force("/s298_fc_tb/uut/G136", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G136", 0);
signal_force("/s298_fc_tb/uut/G136", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G136", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I442 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I442;"));
signal_force("/s298_fc_tb/uut/I442", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I442", 0);
signal_force("/s298_fc_tb/uut/I442", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I442", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G331 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G331;"));
signal_force("/s298_fc_tb/uut/G331", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G331", 0);
signal_force("/s298_fc_tb/uut/G331", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G331", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G88 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G88;"));
signal_force("/s298_fc_tb/uut/G88", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G88", 0);
signal_force("/s298_fc_tb/uut/G88", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G88", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I414 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I414;"));
signal_force("/s298_fc_tb/uut/I414", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I414", 0);
signal_force("/s298_fc_tb/uut/I414", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I414", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G178 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G178;"));
signal_force("/s298_fc_tb/uut/G178", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G178", 0);
signal_force("/s298_fc_tb/uut/G178", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G178", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I449 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I449;"));
signal_force("/s298_fc_tb/uut/I449", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I449", 0);
signal_force("/s298_fc_tb/uut/I449", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I449", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G179 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G179;"));
signal_force("/s298_fc_tb/uut/G179", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G179", 0);
signal_force("/s298_fc_tb/uut/G179", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G179", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I452 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I452;"));
signal_force("/s298_fc_tb/uut/I452", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I452", 0);
signal_force("/s298_fc_tb/uut/I452", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I452", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G357 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G357;"));
signal_force("/s298_fc_tb/uut/G357", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G357", 0);
signal_force("/s298_fc_tb/uut/G357", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G357", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G358 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G358;"));
signal_force("/s298_fc_tb/uut/G358", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G358", 0);
signal_force("/s298_fc_tb/uut/G358", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G358", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G112 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G112;"));
signal_force("/s298_fc_tb/uut/G112", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G112", 0);
signal_force("/s298_fc_tb/uut/G112", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G112", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G335 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G335;"));
signal_force("/s298_fc_tb/uut/G335", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G335", 0);
signal_force("/s298_fc_tb/uut/G335", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G335", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I460 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I460;"));
signal_force("/s298_fc_tb/uut/I460", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I460", 0);
signal_force("/s298_fc_tb/uut/I460", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I460", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G190 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G190;"));
signal_force("/s298_fc_tb/uut/G190", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G190", 0);
signal_force("/s298_fc_tb/uut/G190", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G190", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I463 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I463;"));
signal_force("/s298_fc_tb/uut/I463", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I463", 0);
signal_force("/s298_fc_tb/uut/I463", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I463", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G336 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G336;"));
signal_force("/s298_fc_tb/uut/G336", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G336", 0);
signal_force("/s298_fc_tb/uut/G336", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G336", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G306 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G306;"));
signal_force("/s298_fc_tb/uut/G306", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G306", 0);
signal_force("/s298_fc_tb/uut/G306", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G306", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I466 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I466;"));
signal_force("/s298_fc_tb/uut/I466", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I466", 0);
signal_force("/s298_fc_tb/uut/I466", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I466", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G158 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G158;"));
signal_force("/s298_fc_tb/uut/G158", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G158", 0);
signal_force("/s298_fc_tb/uut/G158", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G158", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I469 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I469;"));
signal_force("/s298_fc_tb/uut/I469", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I469", 0);
signal_force("/s298_fc_tb/uut/I469", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I469", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G307 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G307;"));
signal_force("/s298_fc_tb/uut/G307", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G307", 0);
signal_force("/s298_fc_tb/uut/G307", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G307", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I472 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I472;"));
signal_force("/s298_fc_tb/uut/I472", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I472", 0);
signal_force("/s298_fc_tb/uut/I472", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I472", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G377 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G377;"));
signal_force("/s298_fc_tb/uut/G377", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G377", 0);
signal_force("/s298_fc_tb/uut/G377", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G377", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I476 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I476;"));
signal_force("/s298_fc_tb/uut/I476", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I476", 0);
signal_force("/s298_fc_tb/uut/I476", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I476", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G378 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G378;"));
signal_force("/s298_fc_tb/uut/G378", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G378", 0);
signal_force("/s298_fc_tb/uut/G378", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G378", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G99 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G99;"));
signal_force("/s298_fc_tb/uut/G99", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G99", 0);
signal_force("/s298_fc_tb/uut/G99", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G99", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G395 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G395;"));
signal_force("/s298_fc_tb/uut/G395", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G395", 0);
signal_force("/s298_fc_tb/uut/G395", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G395", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G105 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G105;"));
signal_force("/s298_fc_tb/uut/G105", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G105", 0);
signal_force("/s298_fc_tb/uut/G105", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G105", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G277 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G277;"));
signal_force("/s298_fc_tb/uut/G277", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G277", 0);
signal_force("/s298_fc_tb/uut/G277", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G277", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II272 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II272;"));
signal_force("/s298_fc_tb/uut/II272", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II272", 0);
signal_force("/s298_fc_tb/uut/II272", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II272", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G276 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G276;"));
signal_force("/s298_fc_tb/uut/G276", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G276", 0);
signal_force("/s298_fc_tb/uut/G276", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G276", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I265 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I265;"));
signal_force("/s298_fc_tb/uut/I265", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I265", 0);
signal_force("/s298_fc_tb/uut/I265", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I265", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G284 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G284;"));
signal_force("/s298_fc_tb/uut/G284", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G284", 0);
signal_force("/s298_fc_tb/uut/G284", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G284", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I320 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I320;"));
signal_force("/s298_fc_tb/uut/I320", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I320", 0);
signal_force("/s298_fc_tb/uut/I320", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I320", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G279 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G279;"));
signal_force("/s298_fc_tb/uut/G279", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G279", 0);
signal_force("/s298_fc_tb/uut/G279", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G279", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I285 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I285;"));
signal_force("/s298_fc_tb/uut/I285", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I285", 0);
signal_force("/s298_fc_tb/uut/I285", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I285", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G280 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G280;"));
signal_force("/s298_fc_tb/uut/G280", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G280", 0);
signal_force("/s298_fc_tb/uut/G280", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G280", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I292 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I292;"));
signal_force("/s298_fc_tb/uut/I292", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I292", 0);
signal_force("/s298_fc_tb/uut/I292", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I292", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I322 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I322;"));
signal_force("/s298_fc_tb/uut/I322", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I322", 0);
signal_force("/s298_fc_tb/uut/I322", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I322", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II287 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II287;"));
signal_force("/s298_fc_tb/uut/II287", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II287", 0);
signal_force("/s298_fc_tb/uut/II287", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II287", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I294 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I294;"));
signal_force("/s298_fc_tb/uut/I294", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I294", 0);
signal_force("/s298_fc_tb/uut/I294", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I294", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G134 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G134;"));
signal_force("/s298_fc_tb/uut/G134", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G134", 0);
signal_force("/s298_fc_tb/uut/G134", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G134", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I517 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I517;"));
signal_force("/s298_fc_tb/uut/I517", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I517", 0);
signal_force("/s298_fc_tb/uut/I517", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I517", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G327 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G327;"));
signal_force("/s298_fc_tb/uut/G327", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G327", 0);
signal_force("/s298_fc_tb/uut/G327", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G327", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G86 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G86;"));
signal_force("/s298_fc_tb/uut/G86", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G86", 0);
signal_force("/s298_fc_tb/uut/G86", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G86", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I398 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I398;"));
signal_force("/s298_fc_tb/uut/I398", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I398", 0);
signal_force("/s298_fc_tb/uut/I398", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I398", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G168 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G168;"));
signal_force("/s298_fc_tb/uut/G168", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G168", 0);
signal_force("/s298_fc_tb/uut/G168", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G168", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I524 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I524;"));
signal_force("/s298_fc_tb/uut/I524", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I524", 0);
signal_force("/s298_fc_tb/uut/I524", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I524", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G169 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G169;"));
signal_force("/s298_fc_tb/uut/G169", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G169", 0);
signal_force("/s298_fc_tb/uut/G169", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G169", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I527 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I527;"));
signal_force("/s298_fc_tb/uut/I527", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I527", 0);
signal_force("/s298_fc_tb/uut/I527", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I527", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G353 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G353;"));
signal_force("/s298_fc_tb/uut/G353", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G353", 0);
signal_force("/s298_fc_tb/uut/G353", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G353", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G354 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G354;"));
signal_force("/s298_fc_tb/uut/G354", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G354", 0);
signal_force("/s298_fc_tb/uut/G354", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G354", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G120 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G120;"));
signal_force("/s298_fc_tb/uut/G120", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G120", 0);
signal_force("/s298_fc_tb/uut/G120", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G120", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G347 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G347;"));
signal_force("/s298_fc_tb/uut/G347", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G347", 0);
signal_force("/s298_fc_tb/uut/G347", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G347", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I535 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I535;"));
signal_force("/s298_fc_tb/uut/I535", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I535", 0);
signal_force("/s298_fc_tb/uut/I535", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I535", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G206 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G206;"));
signal_force("/s298_fc_tb/uut/G206", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G206", 0);
signal_force("/s298_fc_tb/uut/G206", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G206", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I538 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I538;"));
signal_force("/s298_fc_tb/uut/I538", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I538", 0);
signal_force("/s298_fc_tb/uut/I538", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I538", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G348 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G348;"));
signal_force("/s298_fc_tb/uut/G348", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G348", 0);
signal_force("/s298_fc_tb/uut/G348", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G348", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G300 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G300;"));
signal_force("/s298_fc_tb/uut/G300", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G300", 0);
signal_force("/s298_fc_tb/uut/G300", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G300", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I541 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I541;"));
signal_force("/s298_fc_tb/uut/I541", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I541", 0);
signal_force("/s298_fc_tb/uut/I541", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I541", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G150 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G150;"));
signal_force("/s298_fc_tb/uut/G150", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G150", 0);
signal_force("/s298_fc_tb/uut/G150", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G150", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I544 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I544;"));
signal_force("/s298_fc_tb/uut/I544", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I544", 0);
signal_force("/s298_fc_tb/uut/I544", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I544", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G301 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G301;"));
signal_force("/s298_fc_tb/uut/G301", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G301", 0);
signal_force("/s298_fc_tb/uut/G301", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G301", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I547 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I547;"));
signal_force("/s298_fc_tb/uut/I547", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I547", 0);
signal_force("/s298_fc_tb/uut/I547", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I547", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G369 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G369;"));
signal_force("/s298_fc_tb/uut/G369", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G369", 0);
signal_force("/s298_fc_tb/uut/G369", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G369", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I551 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I551;"));
signal_force("/s298_fc_tb/uut/I551", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I551", 0);
signal_force("/s298_fc_tb/uut/I551", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I551", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G370 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G370;"));
signal_force("/s298_fc_tb/uut/G370", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G370", 0);
signal_force("/s298_fc_tb/uut/G370", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G370", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G95 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G95;"));
signal_force("/s298_fc_tb/uut/G95", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G95", 0);
signal_force("/s298_fc_tb/uut/G95", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G95", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G391 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G391;"));
signal_force("/s298_fc_tb/uut/G391", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G391", 0);
signal_force("/s298_fc_tb/uut/G391", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G391", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G103 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G103;"));
signal_force("/s298_fc_tb/uut/G103", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G103", 0);
signal_force("/s298_fc_tb/uut/G103", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G103", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G271 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G271;"));
signal_force("/s298_fc_tb/uut/G271", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G271", 0);
signal_force("/s298_fc_tb/uut/G271", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G271", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I230 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I230;"));
signal_force("/s298_fc_tb/uut/I230", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I230", 0);
signal_force("/s298_fc_tb/uut/I230", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I230", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G275 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G275;"));
signal_force("/s298_fc_tb/uut/G275", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G275", 0);
signal_force("/s298_fc_tb/uut/G275", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G275", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I258 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I258;"));
signal_force("/s298_fc_tb/uut/I258", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I258", 0);
signal_force("/s298_fc_tb/uut/I258", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I258", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G288 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G288;"));
signal_force("/s298_fc_tb/uut/G288", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G288", 0);
signal_force("/s298_fc_tb/uut/G288", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G288", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I348 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I348;"));
signal_force("/s298_fc_tb/uut/I348", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I348", 0);
signal_force("/s298_fc_tb/uut/I348", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I348", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G287 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G287;"));
signal_force("/s298_fc_tb/uut/G287", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G287", 0);
signal_force("/s298_fc_tb/uut/G287", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G287", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II341 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II341;"));
signal_force("/s298_fc_tb/uut/II341", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II341", 0);
signal_force("/s298_fc_tb/uut/II341", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II341", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G270 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G270;"));
signal_force("/s298_fc_tb/uut/G270", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G270", 0);
signal_force("/s298_fc_tb/uut/G270", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G270", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I222 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I222;"));
signal_force("/s298_fc_tb/uut/I222", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I222", 0);
signal_force("/s298_fc_tb/uut/I222", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I222", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I350 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I350;"));
signal_force("/s298_fc_tb/uut/I350", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I350", 0);
signal_force("/s298_fc_tb/uut/I350", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I350", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I343 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I343;"));
signal_force("/s298_fc_tb/uut/I343", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I343", 0);
signal_force("/s298_fc_tb/uut/I343", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I343", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G272 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G272;"));
signal_force("/s298_fc_tb/uut/G272", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G272", 0);
signal_force("/s298_fc_tb/uut/G272", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G272", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I237 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I237;"));
signal_force("/s298_fc_tb/uut/I237", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I237", 0);
signal_force("/s298_fc_tb/uut/I237", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I237", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G273 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G273;"));
signal_force("/s298_fc_tb/uut/G273", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G273", 0);
signal_force("/s298_fc_tb/uut/G273", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G273", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I244 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I244;"));
signal_force("/s298_fc_tb/uut/I244", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I244", 0);
signal_force("/s298_fc_tb/uut/I244", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I244", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G274 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G274;"));
signal_force("/s298_fc_tb/uut/G274", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G274", 0);
signal_force("/s298_fc_tb/uut/G274", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G274", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I251 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I251;"));
signal_force("/s298_fc_tb/uut/I251", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I251", 0);
signal_force("/s298_fc_tb/uut/I251", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I251", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I224 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I224;"));
signal_force("/s298_fc_tb/uut/I224", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I224", 0);
signal_force("/s298_fc_tb/uut/I224", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I224", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G124 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G124;"));
signal_force("/s298_fc_tb/uut/G124", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G124", 0);
signal_force("/s298_fc_tb/uut/G124", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G124", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I608 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I608;"));
signal_force("/s298_fc_tb/uut/I608", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I608", 0);
signal_force("/s298_fc_tb/uut/I608", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I608", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G298 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G298;"));
signal_force("/s298_fc_tb/uut/G298", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G298", 0);
signal_force("/s298_fc_tb/uut/G298", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G298", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G231 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G231;"));
signal_force("/s298_fc_tb/uut/G231", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G231", 0);
signal_force("/s298_fc_tb/uut/G231", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G231", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G232 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G232;"));
signal_force("/s298_fc_tb/uut/G232", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G232", 0);
signal_force("/s298_fc_tb/uut/G232", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G232", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G233 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G233;"));
signal_force("/s298_fc_tb/uut/G233", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G233", 0);
signal_force("/s298_fc_tb/uut/G233", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G233", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G234 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G234;"));
signal_force("/s298_fc_tb/uut/G234", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G234", 0);
signal_force("/s298_fc_tb/uut/G234", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G234", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G247 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G247;"));
signal_force("/s298_fc_tb/uut/G247", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G247", 0);
signal_force("/s298_fc_tb/uut/G247", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G247", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G248 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G248;"));
signal_force("/s298_fc_tb/uut/G248", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G248", 0);
signal_force("/s298_fc_tb/uut/G248", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G248", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G263 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G263;"));
signal_force("/s298_fc_tb/uut/G263", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G263", 0);
signal_force("/s298_fc_tb/uut/G263", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G263", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G264 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G264;"));
signal_force("/s298_fc_tb/uut/G264", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G264", 0);
signal_force("/s298_fc_tb/uut/G264", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G264", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G33 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G33;"));
signal_force("/s298_fc_tb/uut/G33", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G33", 0);
signal_force("/s298_fc_tb/uut/G33", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G33", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G107 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G107;"));
signal_force("/s298_fc_tb/uut/G107", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G107", 0);
signal_force("/s298_fc_tb/uut/G107", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G107", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G83 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G83;"));
signal_force("/s298_fc_tb/uut/G83", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G83", 0);
signal_force("/s298_fc_tb/uut/G83", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G83", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G84 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G84;"));
signal_force("/s298_fc_tb/uut/G84", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G84", 0);
signal_force("/s298_fc_tb/uut/G84", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G84", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G85 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G85;"));
signal_force("/s298_fc_tb/uut/G85", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G85", 0);
signal_force("/s298_fc_tb/uut/G85", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G85", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G92 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G92;"));
signal_force("/s298_fc_tb/uut/G92", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G92", 0);
signal_force("/s298_fc_tb/uut/G92", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G92", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G23 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G23;"));
signal_force("/s298_fc_tb/uut/G23", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G23", 0);
signal_force("/s298_fc_tb/uut/G23", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G23", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G214 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G214;"));
signal_force("/s298_fc_tb/uut/G214", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G214", 0);
signal_force("/s298_fc_tb/uut/G214", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G214", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G210 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G210;"));
signal_force("/s298_fc_tb/uut/G210", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G210", 0);
signal_force("/s298_fc_tb/uut/G210", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G210", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G17 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G17;"));
signal_force("/s298_fc_tb/uut/G17", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G17", 0);
signal_force("/s298_fc_tb/uut/G17", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G17", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G15 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G15;"));
signal_force("/s298_fc_tb/uut/G15", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G15", 0);
signal_force("/s298_fc_tb/uut/G15", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G15", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G240 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G240;"));
signal_force("/s298_fc_tb/uut/G240", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G240", 0);
signal_force("/s298_fc_tb/uut/G240", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G240", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G266 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G266;"));
signal_force("/s298_fc_tb/uut/G266", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G266", 0);
signal_force("/s298_fc_tb/uut/G266", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G266", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G229 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G229;"));
signal_force("/s298_fc_tb/uut/G229", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G229", 0);
signal_force("/s298_fc_tb/uut/G229", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G229", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G245 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G245;"));
signal_force("/s298_fc_tb/uut/G245", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G245", 0);
signal_force("/s298_fc_tb/uut/G245", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G245", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G253 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G253;"));
signal_force("/s298_fc_tb/uut/G253", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G253", 0);
signal_force("/s298_fc_tb/uut/G253", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G253", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I533 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I533;"));
signal_force("/s298_fc_tb/uut/I533", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I533", 0);
signal_force("/s298_fc_tb/uut/I533", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I533", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G227 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G227;"));
signal_force("/s298_fc_tb/uut/G227", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G227", 0);
signal_force("/s298_fc_tb/uut/G227", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G227", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G243 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G243;"));
signal_force("/s298_fc_tb/uut/G243", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G243", 0);
signal_force("/s298_fc_tb/uut/G243", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G243", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G249 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G249;"));
signal_force("/s298_fc_tb/uut/G249", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G249", 0);
signal_force("/s298_fc_tb/uut/G249", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G249", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G265 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G265;"));
signal_force("/s298_fc_tb/uut/G265", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G265", 0);
signal_force("/s298_fc_tb/uut/G265", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G265", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G236 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G236;"));
signal_force("/s298_fc_tb/uut/G236", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G236", 0);
signal_force("/s298_fc_tb/uut/G236", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G236", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G237 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G237;"));
signal_force("/s298_fc_tb/uut/G237", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G237", 0);
signal_force("/s298_fc_tb/uut/G237", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G237", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G252 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G252;"));
signal_force("/s298_fc_tb/uut/G252", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G252", 0);
signal_force("/s298_fc_tb/uut/G252", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G252", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II527 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II527;"));
signal_force("/s298_fc_tb/uut/II527", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II527", 0);
signal_force("/s298_fc_tb/uut/II527", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II527", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G212 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G212;"));
signal_force("/s298_fc_tb/uut/G212", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G212", 0);
signal_force("/s298_fc_tb/uut/G212", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G212", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G16 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G16;"));
signal_force("/s298_fc_tb/uut/G16", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G16", 0);
signal_force("/s298_fc_tb/uut/G16", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G16", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G251 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G251;"));
signal_force("/s298_fc_tb/uut/G251", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G251", 0);
signal_force("/s298_fc_tb/uut/G251", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G251", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I512 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I512;"));
signal_force("/s298_fc_tb/uut/I512", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I512", 0);
signal_force("/s298_fc_tb/uut/I512", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I512", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II538 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II538;"));
signal_force("/s298_fc_tb/uut/II538", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II538", 0);
signal_force("/s298_fc_tb/uut/II538", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II538", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G228 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G228;"));
signal_force("/s298_fc_tb/uut/G228", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G228", 0);
signal_force("/s298_fc_tb/uut/G228", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G228", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G244 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G244;"));
signal_force("/s298_fc_tb/uut/G244", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G244", 0);
signal_force("/s298_fc_tb/uut/G244", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G244", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G256 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G256;"));
signal_force("/s298_fc_tb/uut/G256", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G256", 0);
signal_force("/s298_fc_tb/uut/G256", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G256", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G230 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G230;"));
signal_force("/s298_fc_tb/uut/G230", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G230", 0);
signal_force("/s298_fc_tb/uut/G230", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G230", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G235 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G235;"));
signal_force("/s298_fc_tb/uut/G235", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G235", 0);
signal_force("/s298_fc_tb/uut/G235", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G235", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G246 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G246;"));
signal_force("/s298_fc_tb/uut/G246", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G246", 0);
signal_force("/s298_fc_tb/uut/G246", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G246", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I515 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I515;"));
signal_force("/s298_fc_tb/uut/I515", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I515", 0);
signal_force("/s298_fc_tb/uut/I515", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I515", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G261 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G261;"));
signal_force("/s298_fc_tb/uut/G261", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G261", 0);
signal_force("/s298_fc_tb/uut/G261", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G261", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G208 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G208;"));
signal_force("/s298_fc_tb/uut/G208", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G208", 0);
signal_force("/s298_fc_tb/uut/G208", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G208", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G14 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G14;"));
signal_force("/s298_fc_tb/uut/G14", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G14", 0);
signal_force("/s298_fc_tb/uut/G14", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G14", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I495 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I495;"));
signal_force("/s298_fc_tb/uut/I495", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I495", 0);
signal_force("/s298_fc_tb/uut/I495", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I495", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G255 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G255;"));
signal_force("/s298_fc_tb/uut/G255", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G255", 0);
signal_force("/s298_fc_tb/uut/G255", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G255", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G257 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G257;"));
signal_force("/s298_fc_tb/uut/G257", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G257", 0);
signal_force("/s298_fc_tb/uut/G257", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G257", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I537 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I537;"));
signal_force("/s298_fc_tb/uut/I537", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I537", 0);
signal_force("/s298_fc_tb/uut/I537", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I537", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G226 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G226;"));
signal_force("/s298_fc_tb/uut/G226", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G226", 0);
signal_force("/s298_fc_tb/uut/G226", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G226", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G242 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G242;"));
signal_force("/s298_fc_tb/uut/G242", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G242", 0);
signal_force("/s298_fc_tb/uut/G242", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G242", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I553 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I553;"));
signal_force("/s298_fc_tb/uut/I553", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I553", 0);
signal_force("/s298_fc_tb/uut/I553", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I553", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G241 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G241;"));
signal_force("/s298_fc_tb/uut/G241", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G241", 0);
signal_force("/s298_fc_tb/uut/G241", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G241", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G267 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G267;"));
signal_force("/s298_fc_tb/uut/G267", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G267", 0);
signal_force("/s298_fc_tb/uut/G267", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G267", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G238 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G238;"));
signal_force("/s298_fc_tb/uut/G238", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G238", 0);
signal_force("/s298_fc_tb/uut/G238", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G238", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G239 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G239;"));
signal_force("/s298_fc_tb/uut/G239", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G239", 0);
signal_force("/s298_fc_tb/uut/G239", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G239", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G254 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G254;"));
signal_force("/s298_fc_tb/uut/G254", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G254", 0);
signal_force("/s298_fc_tb/uut/G254", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G254", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I518 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I518;"));
signal_force("/s298_fc_tb/uut/I518", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I518", 0);
signal_force("/s298_fc_tb/uut/I518", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I518", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I521 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I521;"));
signal_force("/s298_fc_tb/uut/I521", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I521", 0);
signal_force("/s298_fc_tb/uut/I521", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I521", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II524 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II524;"));
signal_force("/s298_fc_tb/uut/II524", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II524", 0);
signal_force("/s298_fc_tb/uut/II524", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II524", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G258 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G258;"));
signal_force("/s298_fc_tb/uut/G258", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G258", 0);
signal_force("/s298_fc_tb/uut/G258", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G258", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G259 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G259;"));
signal_force("/s298_fc_tb/uut/G259", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G259", 0);
signal_force("/s298_fc_tb/uut/G259", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G259", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G260 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G260;"));
signal_force("/s298_fc_tb/uut/G260", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G260", 0);
signal_force("/s298_fc_tb/uut/G260", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G260", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal G26 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("G26;"));
signal_force("/s298_fc_tb/uut/G26", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/G26", 0);
signal_force("/s298_fc_tb/uut/G26", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/G26", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I546 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I546;"));
signal_force("/s298_fc_tb/uut/I546", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I546", 0);
signal_force("/s298_fc_tb/uut/I546", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I546", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I300 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I300;"));
signal_force("/s298_fc_tb/uut/I300", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I300", 0);
signal_force("/s298_fc_tb/uut/I300", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I300", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I314 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I314;"));
signal_force("/s298_fc_tb/uut/I314", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I314", 0);
signal_force("/s298_fc_tb/uut/I314", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I314", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I307 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I307;"));
signal_force("/s298_fc_tb/uut/I307", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I307", 0);
signal_force("/s298_fc_tb/uut/I307", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I307", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II335 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II335;"));
signal_force("/s298_fc_tb/uut/II335", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II335", 0);
signal_force("/s298_fc_tb/uut/II335", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II335", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I328 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I328;"));
signal_force("/s298_fc_tb/uut/I328", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I328", 0);
signal_force("/s298_fc_tb/uut/I328", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I328", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I209 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I209;"));
signal_force("/s298_fc_tb/uut/I209", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I209", 0);
signal_force("/s298_fc_tb/uut/I209", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I209", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal II321 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("II321;"));
signal_force("/s298_fc_tb/uut/II321", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/II321", 0);
signal_force("/s298_fc_tb/uut/II321", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/II321", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I286 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I286;"));
signal_force("/s298_fc_tb/uut/I286", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I286", 0);
signal_force("/s298_fc_tb/uut/I286", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I286", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I293 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I293;"));
signal_force("/s298_fc_tb/uut/I293", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I293", 0);
signal_force("/s298_fc_tb/uut/I293", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I293", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I349 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I349;"));
signal_force("/s298_fc_tb/uut/I349", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I349", 0);
signal_force("/s298_fc_tb/uut/I349", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I349", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I342 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I342;"));
signal_force("/s298_fc_tb/uut/I342", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I342", 0);
signal_force("/s298_fc_tb/uut/I342", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I342", 0);
writeline(out_file, s_a_line);
--------------------------------------------------------------------------------
-- Testing signal I223 with stuck-at-1 and stuck-at-0
write(s_a_line,string'("I223;"));
signal_force("/s298_fc_tb/uut/I223", "1", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
write(s_a_line,string'(";"));
wait for clock_period;
signal_release("/s298_fc_tb/uut/I223", 0);
signal_force("/s298_fc_tb/uut/I223", "0", open, freeze, open, 0);
BIST_start_in <= '1';
wait for clock_period;
BIST_start_in <= '0';
wait until BIST_Done_out = '1';
wait for 0.2*clock_period;
write(s_a_line, NOT BIST_result_out);
wait for clock_period;
signal_release("/s298_fc_tb/uut/I223", 0);
writeline(out_file, s_a_line);
