------------------------------------------------------------------------
--#LIS#
--Author: Sebastian Kroesche
--Date: 20.1.2016 
--Description: Implementation of ISCAS89 s1196 circuit with
--             D-type flip-flops
--             generated with bench2vhdl
--Circuit statistics
--# 14 inputs
--# 14 outputs
--# 18 D-type flipflops
--# 141 inverters
--# 388 gates (118 ANDs + 119 NANDs + 101 ORs + 50 NORs)
------------------------------------------------------------------------
library IEEE;
 use IEEE.std_logic_1164.all; 
 
library lis_lib;
 use lis_lib.ser_bist.all; 
 
entity s1196 is
port (
clk : in std_logic; 
reset : in std_logic; 
G0: in std_logic; 
G1: in std_logic; 
G2: in std_logic; 
G3: in std_logic; 
G4: in std_logic; 
G5: in std_logic; 
G6: in std_logic; 
G7: in std_logic; 
G8: in std_logic; 
G9: in std_logic; 
G10: in std_logic; 
G11: in std_logic; 
G12: in std_logic; 
G13: in std_logic; 
G546: out std_logic; 
G539: out std_logic; 
G550: out std_logic; 
G551: out std_logic; 
G552: out std_logic; 
G547: out std_logic; 
G548: out std_logic; 
G549: out std_logic; 
G530: out std_logic; 
G45: out std_logic; 
G542: out std_logic; 
G532: out std_logic; 
G535: out std_logic; 
G537: out std_logic 
);
end entity; 

architecture rtl of s1196 is
begin

--Flip-flops (total number: 18)
DFF_0:	 lis_dff port map( clk => clk, Q_out => G29, D_in => G502, reset => reset );
DFF_1:	 lis_dff port map( clk => clk, Q_out => G30, D_in => G503, reset => reset );
DFF_2:	 lis_dff port map( clk => clk, Q_out => G31, D_in => G504, reset => reset );
DFF_3:	 lis_dff port map( clk => clk, Q_out => G32, D_in => G505, reset => reset );
DFF_4:	 lis_dff port map( clk => clk, Q_out => G33, D_in => G506, reset => reset );
DFF_5:	 lis_dff port map( clk => clk, Q_out => G34, D_in => G507, reset => reset );
DFF_6:	 lis_dff port map( clk => clk, Q_out => G35, D_in => G508, reset => reset );
DFF_7:	 lis_dff port map( clk => clk, Q_out => G36, D_in => G509, reset => reset );
DFF_8:	 lis_dff port map( clk => clk, Q_out => G37, D_in => G510, reset => reset );
DFF_9:	 lis_dff port map( clk => clk, Q_out => G38, D_in => G511, reset => reset );
DFF_10:	 lis_dff port map( clk => clk, Q_out => G39, D_in => G512, reset => reset );
DFF_11:	 lis_dff port map( clk => clk, Q_out => G40, D_in => G513, reset => reset );
DFF_12:	 lis_dff port map( clk => clk, Q_out => G41, D_in => G514, reset => reset );
DFF_13:	 lis_dff port map( clk => clk, Q_out => G42, D_in => G515, reset => reset );
DFF_14:	 lis_dff port map( clk => clk, Q_out => G43, D_in => G516, reset => reset );
DFF_15:	 lis_dff port map( clk => clk, Q_out => G44, D_in => G517, reset => reset );
DFF_16:	 lis_dff port map( clk => clk, Q_out => G45, D_in => G518, reset => reset );
DFF_17:	 lis_dff port map( clk => clk, Q_out => G46, D_in => G519, reset => reset );

--Inverters (total number: 141)
INV_0:	 lis_not port map( A => G0, Z => G520 );
INV_1:	 lis_not port map( A => G1, Z => G521 );
INV_2:	 lis_not port map( A => G2, Z => G522 );
INV_3:	 lis_not port map( A => G3, Z => G524 );
INV_4:	 lis_not port map( A => G4, Z => I156 );
INV_5:	 lis_not port map( A => I156, Z => G334 );
INV_6:	 lis_not port map( A => G4, Z => G527 );
INV_7:	 lis_not port map( A => G5, Z => G528 );
INV_8:	 lis_not port map( A => G6, Z => G529 );
INV_9:	 lis_not port map( A => G7, Z => G531 );
INV_10:	 lis_not port map( A => G8, Z => G533 );
INV_11:	 lis_not port map( A => G9, Z => G536 );
INV_12:	 lis_not port map( A => G10, Z => G538 );
INV_13:	 lis_not port map( A => G11, Z => G540 );
INV_14:	 lis_not port map( A => G12, Z => G541 );
INV_15:	 lis_not port map( A => G13, Z => G543 );
INV_16:	 lis_not port map( A => G30, Z => G476 );
INV_17:	 lis_not port map( A => G30, Z => G484 );
INV_18:	 lis_not port map( A => G40, Z => G125 );
INV_19:	 lis_not port map( A => G33, Z => G140 );
INV_20:	 lis_not port map( A => G41, Z => G546 );
INV_21:	 lis_not port map( A => G42, Z => G132 );
INV_22:	 lis_not port map( A => G43, Z => G70 );
INV_23:	 lis_not port map( A => G44, Z => G67 );
INV_24:	 lis_not port map( A => G29, Z => G99 );
INV_25:	 lis_not port map( A => G57, Z => G475 );
INV_26:	 lis_not port map( A => G58, Z => G59 );
INV_27:	 lis_not port map( A => G524, Z => G228 );
INV_28:	 lis_not port map( A => G271, Z => G272 );
INV_29:	 lis_not port map( A => G97, Z => G98 );
INV_30:	 lis_not port map( A => G134, Z => G135 );
INV_31:	 lis_not port map( A => G528, Z => I218 );
INV_32:	 lis_not port map( A => I218, Z => G333 );
INV_33:	 lis_not port map( A => G54, Z => G55 );
INV_34:	 lis_not port map( A => G529, Z => G165 );
INV_35:	 lis_not port map( A => G71, Z => G72 );
INV_36:	 lis_not port map( A => G274, Z => G236 );
INV_37:	 lis_not port map( A => G274, Z => G275 );
INV_38:	 lis_not port map( A => G538, Z => I249 );
INV_39:	 lis_not port map( A => I249, Z => G370 );
INV_40:	 lis_not port map( A => G74, Z => G75 );
INV_41:	 lis_not port map( A => G190, Z => G490 );
INV_42:	 lis_not port map( A => G241, Z => G482 );
INV_43:	 lis_not port map( A => G522, Z => G153 );
INV_44:	 lis_not port map( A => G193, Z => G192 );
INV_45:	 lis_not port map( A => G122, Z => G123 );
INV_46:	 lis_not port map( A => G209, Z => I272 );
INV_47:	 lis_not port map( A => I272, Z => G458 );
INV_48:	 lis_not port map( A => G238, Z => I276 );
INV_49:	 lis_not port map( A => I276, Z => G332 );
INV_50:	 lis_not port map( A => G272, Z => I280 );
INV_51:	 lis_not port map( A => I280, Z => G309 );
INV_52:	 lis_not port map( A => G135, Z => I287 );
INV_53:	 lis_not port map( A => I287, Z => G347 );
INV_54:	 lis_not port map( A => G195, Z => G498 );
INV_55:	 lis_not port map( A => G77, Z => G78 );
INV_56:	 lis_not port map( A => G198, Z => I295 );
INV_57:	 lis_not port map( A => I295, Z => G459 );
INV_58:	 lis_not port map( A => G200, Z => G199 );
INV_59:	 lis_not port map( A => G89, Z => G90 );
INV_60:	 lis_not port map( A => G222, Z => G221 );
INV_61:	 lis_not port map( A => G224, Z => G223 );
INV_62:	 lis_not port map( A => G239, Z => I316 );
INV_63:	 lis_not port map( A => I316, Z => G369 );
INV_64:	 lis_not port map( A => G235, Z => G234 );
INV_65:	 lis_not port map( A => G135, Z => I327 );
INV_66:	 lis_not port map( A => I327, Z => G435 );
INV_67:	 lis_not port map( A => G236, Z => I330 );
INV_68:	 lis_not port map( A => I330, Z => G441 );
INV_69:	 lis_not port map( A => G49, Z => G50 );
INV_70:	 lis_not port map( A => G9, Z => G130 );
INV_71:	 lis_not port map( A => G156, Z => G501 );
INV_72:	 lis_not port map( A => G276, Z => G477 );
INV_73:	 lis_not port map( A => G276, Z => G485 );
INV_74:	 lis_not port map( A => G77, Z => I352 );
INV_75:	 lis_not port map( A => I352, Z => G299 );
INV_76:	 lis_not port map( A => G205, Z => G497 );
INV_77:	 lis_not port map( A => G1, Z => I371 );
INV_78:	 lis_not port map( A => I371, Z => G335 );
INV_79:	 lis_not port map( A => G520, Z => I374 );
INV_80:	 lis_not port map( A => I374, Z => G456 );
INV_81:	 lis_not port map( A => G86, Z => G87 );
INV_82:	 lis_not port map( A => G199, Z => I386 );
INV_83:	 lis_not port map( A => I386, Z => G414 );
INV_84:	 lis_not port map( A => G68, Z => G486 );
INV_85:	 lis_not port map( A => G232, Z => G231 );
INV_86:	 lis_not port map( A => G161, Z => G160 );
INV_87:	 lis_not port map( A => G50, Z => G265 );
INV_88:	 lis_not port map( A => G63, Z => G64 );
INV_89:	 lis_not port map( A => G181, Z => G180 );
INV_90:	 lis_not port map( A => G456, Z => G107 );
INV_91:	 lis_not port map( A => G208, Z => G207 );
INV_92:	 lis_not port map( A => G168, Z => G167 );
INV_93:	 lis_not port map( A => G206, Z => G124 );
INV_94:	 lis_not port map( A => G204, Z => G203 );
INV_95:	 lis_not port map( A => G273, Z => G489 );
INV_96:	 lis_not port map( A => G273, Z => G495 );
INV_97:	 lis_not port map( A => G357, Z => G177 );
INV_98:	 lis_not port map( A => G213, Z => G212 );
INV_99:	 lis_not port map( A => G218, Z => I493 );
INV_100:	 lis_not port map( A => I493, Z => G404 );
INV_101:	 lis_not port map( A => G124, Z => I502 );
INV_102:	 lis_not port map( A => I502, Z => G468 );
INV_103:	 lis_not port map( A => G495, Z => G173 );
INV_104:	 lis_not port map( A => G534, Z => G487 );
INV_105:	 lis_not port map( A => G468, Z => I529 );
INV_106:	 lis_not port map( A => I529, Z => G149 );
INV_107:	 lis_not port map( A => G79, Z => I536 );
INV_108:	 lis_not port map( A => I536, Z => G446 );
INV_109:	 lis_not port map( A => G173, Z => G494 );
INV_110:	 lis_not port map( A => G173, Z => G500 );
INV_111:	 lis_not port map( A => G215, Z => G214 );
INV_112:	 lis_not port map( A => G62, Z => G492 );
INV_113:	 lis_not port map( A => G182, Z => G483 );
INV_114:	 lis_not port map( A => G281, Z => G282 );
INV_115:	 lis_not port map( A => G176, Z => I573 );
INV_116:	 lis_not port map( A => I573, Z => G403 );
INV_117:	 lis_not port map( A => G175, Z => I576 );
INV_118:	 lis_not port map( A => I576, Z => G447 );
INV_119:	 lis_not port map( A => G194, Z => G479 );
INV_120:	 lis_not port map( A => G194, Z => G491 );
INV_121:	 lis_not port map( A => G553, Z => G554 );
INV_122:	 lis_not port map( A => G171, Z => G170 );
INV_123:	 lis_not port map( A => G171, Z => G172 );
INV_124:	 lis_not port map( A => G526, Z => G525 );
INV_125:	 lis_not port map( A => G544, Z => G493 );
INV_126:	 lis_not port map( A => G544, Z => G545 );
INV_127:	 lis_not port map( A => G172, Z => G488 );
INV_128:	 lis_not port map( A => G280, Z => G499 );
INV_129:	 lis_not port map( A => G120, Z => I624 );
INV_130:	 lis_not port map( A => I624, Z => G303 );
INV_131:	 lis_not port map( A => G179, Z => G480 );
INV_132:	 lis_not port map( A => G188, Z => I631 );
INV_133:	 lis_not port map( A => I631, Z => G336 );
INV_134:	 lis_not port map( A => G188, Z => G496 );
INV_135:	 lis_not port map( A => G496, Z => G174 );
INV_136:	 lis_not port map( A => G174, Z => I662 );
INV_137:	 lis_not port map( A => I662, Z => G405 );
INV_138:	 lis_not port map( A => G279, Z => G478 );
INV_139:	 lis_not port map( A => G145, Z => I692 );
INV_140:	 lis_not port map( A => I692, Z => G432 );

--AND-gates (total number: 118)
AND2_0:	 LIS_AND2 port map( A => G6, B => G31, Z => G359);
AND2_1:	 LIS_AND2 port map( A => G163, B => G3, Z => G469);
AND2_2:	 LIS_AND2 port map( A => G529, B => G531, Z => G461);
AND2_3:	 LIS_AND2 port map( A => G524, B => G67, Z => G431);
AND2_4:	 LIS_AND2 port map( A => G129, B => G77, Z => G362);
AND2_5:	 LIS_AND2 port map( A => G288, B => G240, Z => G81);
AND2_6:	 LIS_AND2 port map( A => G97, B => G55, Z => G348);
AND4_0:	 LIS_AND4 port map( A => G8, B => G135, C => G37, D => G164, Z => G352 );
AND2_7:	 LIS_AND2 port map( A => G163, B => G164, Z => G511);
AND2_8:	 LIS_AND2 port map( A => G9, B => G211, Z => G379);
AND3_0:	 LIS_AND3 port map( A => G529, B => G7, C => G49, Z => G385 );
AND2_9:	 LIS_AND2 port map( A => G533, B => G75, Z => G376);
AND3_1:	 LIS_AND3 port map( A => G6, B => G274, C => G75, Z => G387 );
AND2_10:	 LIS_AND2 port map( A => G192, B => G538, Z => G462);
AND2_11:	 LIS_AND2 port map( A => G123, B => G77, Z => G436);
AND2_12:	 LIS_AND2 port map( A => G77, B => G205, Z => G363);
AND2_13:	 LIS_AND2 port map( A => G1, B => G205, Z => G410);
AND2_14:	 LIS_AND2 port map( A => G520, B => G1, Z => G399);
AND2_15:	 LIS_AND2 port map( A => G66, B => G229, Z => G437);
AND2_16:	 LIS_AND2 port map( A => G6, B => G104, Z => G307);
AND2_17:	 LIS_AND2 port map( A => G524, B => G78, Z => G306);
AND2_18:	 LIS_AND2 port map( A => G122, B => G219, Z => G283);
AND3_2:	 LIS_AND3 port map( A => G533, B => G199, C => G209, Z => G339 );
AND3_3:	 LIS_AND3 port map( A => G136, B => G9, C => G190, Z => G472 );
AND4_1:	 LIS_AND4 port map( A => G524, B => G169, C => G221, D => G234, Z => G351 );
AND2_19:	 LIS_AND2 port map( A => G38, B => G234, Z => G440);
AND3_4:	 LIS_AND3 port map( A => G9, B => G100, C => G34, Z => G382 );
AND2_20:	 LIS_AND2 port map( A => G536, B => G85, Z => G386);
AND2_21:	 LIS_AND2 port map( A => G90, B => G50, Z => G321);
AND2_22:	 LIS_AND2 port map( A => G89, B => G50, Z => G378);
AND3_5:	 LIS_AND3 port map( A => G191, B => G103, C => G112, Z => G471 );
AND2_23:	 LIS_AND2 port map( A => G90, B => G56, Z => G377);
AND2_24:	 LIS_AND2 port map( A => G7, B => G83, Z => G358);
AND2_25:	 LIS_AND2 port map( A => G0, B => G277, Z => G400);
AND2_26:	 LIS_AND2 port map( A => G5, B => G151, Z => G308);
AND2_27:	 LIS_AND2 port map( A => G48, B => G59, Z => G411);
AND2_28:	 LIS_AND2 port map( A => G197, B => G201, Z => G413);
AND2_29:	 LIS_AND2 port map( A => G165, B => G231, Z => G434);
AND2_30:	 LIS_AND2 port map( A => G34, B => G160, Z => G373);
AND2_31:	 LIS_AND2 port map( A => G265, B => G232, Z => G357);
AND3_6:	 LIS_AND3 port map( A => G64, B => G78, C => G211, Z => G444 );
AND2_32:	 LIS_AND2 port map( A => G6, B => G202, Z => G361);
AND2_33:	 LIS_AND2 port map( A => G2, B => G82, Z => G346);
AND2_34:	 LIS_AND2 port map( A => G4, B => G107, Z => G457);
AND2_35:	 LIS_AND2 port map( A => G2, B => G109, Z => G364);
AND2_36:	 LIS_AND2 port map( A => G53, B => G225, Z => G445);
AND2_37:	 LIS_AND2 port map( A => G3, B => G207, Z => G412);
AND3_7:	 LIS_AND3 port map( A => G161, B => G168, C => G267, Z => G371 );
AND3_8:	 LIS_AND3 port map( A => G11, B => G92, C => G163, Z => G353 );
AND2_38:	 LIS_AND2 port map( A => G11, B => G114, Z => G388);
AND2_39:	 LIS_AND2 port map( A => G11, B => G143, Z => G473);
AND2_40:	 LIS_AND2 port map( A => G213, B => G257, Z => G331);
AND2_41:	 LIS_AND2 port map( A => G51, B => G225, Z => G429);
AND2_42:	 LIS_AND2 port map( A => G6, B => G93, Z => G380);
AND2_43:	 LIS_AND2 port map( A => G8, B => G106, Z => G360);
AND2_44:	 LIS_AND2 port map( A => G202, B => G203, Z => G338);
AND2_45:	 LIS_AND2 port map( A => G270, B => G167, Z => G337);
AND2_46:	 LIS_AND2 port map( A => G8, B => G270, Z => G340);
AND3_9:	 LIS_AND3 port map( A => G522, B => G105, C => G196, Z => G322 );
AND2_47:	 LIS_AND2 port map( A => G248, B => G249, Z => G330);
AND2_48:	 LIS_AND2 port map( A => G177, B => G196, Z => G430);
AND3_10:	 LIS_AND3 port map( A => G111, B => G189, C => G195, Z => G344 );
AND2_49:	 LIS_AND2 port map( A => G212, B => G227, Z => G428);
AND2_50:	 LIS_AND2 port map( A => G6, B => G108, Z => G349);
AND3_11:	 LIS_AND3 port map( A => G2, B => G81, C => G115, Z => G460 );
AND2_51:	 LIS_AND2 port map( A => G521, B => G148, Z => G463);
AND2_52:	 LIS_AND2 port map( A => G127, B => G34, Z => G393);
AND2_53:	 LIS_AND2 port map( A => G528, B => G149, Z => G470);
AND2_54:	 LIS_AND2 port map( A => G531, B => G118, Z => G341);
AND2_55:	 LIS_AND2 port map( A => G73, B => G197, Z => G342);
AND2_56:	 LIS_AND2 port map( A => G522, B => G183, Z => G324);
AND2_57:	 LIS_AND2 port map( A => G2, B => G144, Z => G323);
AND2_58:	 LIS_AND2 port map( A => G0, B => G214, Z => G354);
AND2_59:	 LIS_AND2 port map( A => G180, B => G182, Z => G312);
AND2_60:	 LIS_AND2 port map( A => G250, B => G251, Z => G315);
AND2_61:	 LIS_AND2 port map( A => G242, B => G77, Z => G474);
AND3_12:	 LIS_AND3 port map( A => G2, B => G528, C => G147, Z => G343 );
AND2_62:	 LIS_AND2 port map( A => G52, B => G158, Z => G304);
AND3_13:	 LIS_AND3 port map( A => G94, B => G156, C => G158, Z => G398 );
AND3_14:	 LIS_AND3 port map( A => G282, B => G137, C => G156, Z => G365 );
AND3_15:	 LIS_AND3 port map( A => G13, B => G282, C => G70, Z => G417 );
AND3_16:	 LIS_AND3 port map( A => G117, B => G135, C => G157, Z => G290 );
AND3_17:	 LIS_AND3 port map( A => G4, B => G39, C => G157, Z => G327 );
AND2_63:	 LIS_AND2 port map( A => G126, B => G157, Z => G367);
AND3_18:	 LIS_AND3 port map( A => G101, B => G98, C => G157, Z => G397 );
AND3_19:	 LIS_AND3 port map( A => G541, B => G554, C => G187, Z => G451 );
AND2_64:	 LIS_AND2 port map( A => G87, B => G172, Z => G406);
AND3_20:	 LIS_AND3 port map( A => G524, B => G60, C => G172, Z => G418 );
AND2_65:	 LIS_AND2 port map( A => G545, B => G186, Z => G453);
AND3_21:	 LIS_AND3 port map( A => G2, B => G119, C => G156, Z => G289 );
AND3_22:	 LIS_AND3 port map( A => G0, B => G178, C => G179, Z => G311 );
AND2_66:	 LIS_AND2 port map( A => G154, B => G183, Z => G402);
AND2_67:	 LIS_AND2 port map( A => G91, B => G154, Z => G433);
AND2_68:	 LIS_AND2 port map( A => G88, B => G154, Z => G449);
AND2_69:	 LIS_AND2 port map( A => G526, B => G184, Z => G452);
AND2_70:	 LIS_AND2 port map( A => G150, B => G156, Z => G329);
AND2_71:	 LIS_AND2 port map( A => G138, B => G155, Z => G291);
AND3_23:	 LIS_AND3 port map( A => G5, B => G102, C => G155, Z => G328 );
AND2_72:	 LIS_AND2 port map( A => G125, B => G155, Z => G366);
AND3_24:	 LIS_AND3 port map( A => G116, B => G275, C => G155, Z => G372 );
AND2_73:	 LIS_AND2 port map( A => G131, B => G155, Z => G383);
AND2_74:	 LIS_AND2 port map( A => G132, B => G155, Z => G392);
AND3_25:	 LIS_AND3 port map( A => G76, B => G272, C => G155, Z => G396 );
AND3_26:	 LIS_AND3 port map( A => G2, B => G110, C => G155, Z => G401 );
AND3_27:	 LIS_AND3 port map( A => G0, B => G80, C => G155, Z => G422 );
AND3_28:	 LIS_AND3 port map( A => G146, B => G142, C => G165, Z => G415 );
AND2_75:	 LIS_AND2 port map( A => G146, B => G176, Z => G425);
AND3_29:	 LIS_AND3 port map( A => G8, B => G146, C => G133, Z => G438 );
AND3_30:	 LIS_AND3 port map( A => G78, B => G174, C => G177, Z => G424 );
AND2_76:	 LIS_AND2 port map( A => G174, B => G175, Z => G439);
AND2_77:	 LIS_AND2 port map( A => G159, B => G245, Z => G317);
AND3_31:	 LIS_AND3 port map( A => G37, B => G162, C => G38, Z => G426 );
AND2_78:	 LIS_AND2 port map( A => G47, B => G162, Z => G443);
AND2_79:	 LIS_AND2 port map( A => G61, B => G167, Z => G416);
AND3_32:	 LIS_AND3 port map( A => G541, B => G95, C => G165, Z => G427 );
AND2_80:	 LIS_AND2 port map( A => G541, B => G121, Z => G442);
AND2_81:	 LIS_AND2 port map( A => G541, B => G128, Z => G423);
AND2_82:	 LIS_AND2 port map( A => G139, B => G153, Z => G448);

--OR-gates (total number: 101)
OR2_0:	 LIS_OR2 port map( A => G3, B => G5, Z => G419 );
OR2_1:	 LIS_OR2 port map( A => G6, B => G30, Z => G193 );
OR2_2:	 LIS_OR2 port map( A => G5, B => G58, Z => G394 );
OR2_3:	 LIS_OR2 port map( A => G6, B => G117, Z => G407 );
OR2_4:	 LIS_OR2 port map( A => G527, B => G57, Z => G314 );
OR2_5:	 LIS_OR2 port map( A => G4, B => G134, Z => G395 );
OR2_6:	 LIS_OR2 port map( A => G1, B => G528, Z => G288 );
OR2_7:	 LIS_OR2 port map( A => G4, B => G529, Z => G302 );
OR2_8:	 LIS_OR2 port map( A => G533, B => G31, Z => G224 );
OR2_9:	 LIS_OR2 port map( A => G11, B => G116, Z => G355 );
OR2_10:	 LIS_OR2 port map( A => G531, B => G536, Z => G316 );
OR2_11:	 LIS_OR2 port map( A => G6, B => G536, Z => G350 );
OR2_12:	 LIS_OR2 port map( A => G533, B => G536, Z => G368 );
OR2_13:	 LIS_OR2 port map( A => G7, B => G71, Z => G381 );
OR2_14:	 LIS_OR2 port map( A => G529, B => G71, Z => G384 );
OR2_15:	 LIS_OR2 port map( A => G9, B => G274, Z => G389 );
OR2_16:	 LIS_OR2 port map( A => G536, B => G538, Z => G374 );
OR2_17:	 LIS_OR2 port map( A => G9, B => G540, Z => G286 );
OR2_18:	 LIS_OR2 port map( A => G7, B => G540, Z => G293 );
OR2_19:	 LIS_OR2 port map( A => G10, B => G540, Z => G375 );
OR2_20:	 LIS_OR2 port map( A => G6, B => G476, Z => G356 );
OR2_21:	 LIS_OR2 port map( A => G521, B => G475, Z => G313 );
OR2_22:	 LIS_OR2 port map( A => G522, B => G59, Z => G420 );
OR3_0:	 LIS_OR3 port map( A => G521, B => G2, C => G228, Z => G421 );
OR2_23:	 LIS_OR2 port map( A => G76, B => G272, Z => G320 );
OR2_24:	 LIS_OR2 port map( A => G522, B => G135, Z => G310 );
OR2_25:	 LIS_OR2 port map( A => G529, B => G77, Z => G408 );
OR2_26:	 LIS_OR2 port map( A => G524, B => G55, Z => G305 );
OR2_27:	 LIS_OR2 port map( A => G528, B => G55, Z => G409 );
OR2_28:	 LIS_OR2 port map( A => G89, B => G484, Z => G296 );
OR3_1:	 LIS_OR3 port map( A => G7, B => G536, C => G222, Z => G325 );
OR2_29:	 LIS_OR2 port map( A => G72, B => G536, Z => G464 );
OR2_30:	 LIS_OR2 port map( A => G74, B => G220, Z => G391 );
OR2_31:	 LIS_OR2 port map( A => G538, B => G75, Z => G292 );
OR2_32:	 LIS_OR2 port map( A => G529, B => G226, Z => G345 );
OR2_33:	 LIS_OR2 port map( A => G524, B => G210, Z => G465 );
OR2_34:	 LIS_OR2 port map( A => G122, B => G77, Z => G454 );
OR2_35:	 LIS_OR2 port map( A => G362, B => G529, Z => G269 );
OR2_36:	 LIS_OR2 port map( A => G522, B => G81, Z => G287 );
OR3_2:	 LIS_OR3 port map( A => G6, B => G8, C => G232, Z => G318 );
OR2_37:	 LIS_OR2 port map( A => G533, B => G232, Z => G326 );
OR2_38:	 LIS_OR2 port map( A => G89, B => G50, Z => G390 );
OR2_39:	 LIS_OR2 port map( A => G5, B => G497, Z => G298 );
OR2_40:	 LIS_OR2 port map( A => G87, B => G97, Z => G300 );
OR2_41:	 LIS_OR2 port map( A => G283, B => G528, Z => G261 );
OR2_42:	 LIS_OR2 port map( A => G122, B => G486, Z => G301 );
OR2_43:	 LIS_OR2 port map( A => G351, B => G352, Z => G92 );
OR2_44:	 LIS_OR2 port map( A => G440, B => G441, Z => G47 );
OR2_45:	 LIS_OR2 port map( A => G385, B => G386, Z => G114 );
OR2_46:	 LIS_OR2 port map( A => G64, B => G274, Z => G297 );
OR3_3:	 LIS_OR3 port map( A => G376, B => G377, C => G378, Z => G93 );
OR2_47:	 LIS_OR2 port map( A => G358, B => G359, Z => G106 );
OR2_48:	 LIS_OR2 port map( A => G399, B => G400, Z => G110 );
OR2_49:	 LIS_OR2 port map( A => G78, B => G206, Z => G455 );
OR3_4:	 LIS_OR3 port map( A => G306, B => G307, C => G308, Z => G152 );
OR2_50:	 LIS_OR2 port map( A => G413, B => G414, Z => G60 );
OR2_51:	 LIS_OR2 port map( A => G434, B => G435, Z => G133 );
OR2_52:	 LIS_OR2 port map( A => G321, B => G273, Z => G105 );
OR2_53:	 LIS_OR2 port map( A => G346, B => G347, Z => G108 );
OR3_5:	 LIS_OR3 port map( A => G457, B => G458, C => G459, Z => G115 );
OR2_54:	 LIS_OR2 port map( A => G363, B => G364, Z => G126 );
OR2_55:	 LIS_OR2 port map( A => G444, B => G445, Z => G79 );
OR2_56:	 LIS_OR2 port map( A => G529, B => G489, Z => G319 );
OR2_57:	 LIS_OR2 port map( A => G379, B => G380, Z => G131 );
OR2_58:	 LIS_OR2 port map( A => G337, B => G338, Z => G118 );
OR2_59:	 LIS_OR2 port map( A => G339, B => G340, Z => G73 );
OR2_60:	 LIS_OR2 port map( A => G430, B => G431, Z => G91 );
OR2_61:	 LIS_OR2 port map( A => G348, B => G349, Z => G137 );
OR2_62:	 LIS_OR2 port map( A => G469, B => G470, Z => G242 );
OR2_63:	 LIS_OR2 port map( A => G341, B => G342, Z => G147 );
OR3_6:	 LIS_OR3 port map( A => G528, B => G272, C => G281, Z => G284 );
OR3_7:	 LIS_OR3 port map( A => G1, B => G117, C => G281, Z => G294 );
OR3_8:	 LIS_OR3 port map( A => G322, B => G323, C => G324, Z => G553 );
OR2_64:	 LIS_OR2 port map( A => G353, B => G354, Z => G141 );
OR2_65:	 LIS_OR2 port map( A => G403, B => G404, Z => G142 );
OR2_66:	 LIS_OR2 port map( A => G446, B => G447, Z => G88 );
OR2_67:	 LIS_OR2 port map( A => G343, B => G344, Z => G544 );
OR2_68:	 LIS_OR2 port map( A => G5, B => G479, Z => G285 );
OR2_69:	 LIS_OR2 port map( A => G122, B => G491, Z => G295 );
OR2_70:	 LIS_OR2 port map( A => G12, B => G171, Z => G450 );
OR2_71:	 LIS_OR2 port map( A => G303, B => G304, Z => G150 );
OR2_72:	 LIS_OR2 port map( A => G336, B => G170, Z => G146 );
OR3_9:	 LIS_OR3 port map( A => G451, B => G452, C => G453, Z => G539 );
OR2_73:	 LIS_OR2 port map( A => G371, B => G159, Z => G244 );
OR4_0:	 LIS_OR4 port map( A => G289, B => G290, C => G291, D => G485, Z => G550 );
OR3_10:	 LIS_OR3 port map( A => G327, B => G328, C => G329, Z => G551 );
OR3_11:	 LIS_OR3 port map( A => G365, B => G366, C => G367, Z => G552 );
OR2_74:	 LIS_OR2 port map( A => G382, B => G383, Z => G547 );
OR2_75:	 LIS_OR2 port map( A => G392, B => G393, Z => G548 );
OR4_1:	 LIS_OR4 port map( A => G396, B => G397, C => G398, D => G477, Z => G549 );
OR2_76:	 LIS_OR2 port map( A => G401, B => G402, Z => G530 );
OR2_77:	 LIS_OR2 port map( A => G405, B => G406, Z => G61 );
OR2_78:	 LIS_OR2 port map( A => G424, B => G425, Z => G95 );
OR2_79:	 LIS_OR2 port map( A => G438, B => G439, Z => G121 );
OR2_80:	 LIS_OR2 port map( A => G317, B => G166, Z => G279 );
OR4_2:	 LIS_OR4 port map( A => G415, B => G416, C => G417, D => G418, Z => G128 );
OR2_81:	 LIS_OR2 port map( A => G426, B => G427, Z => G145 );
OR2_82:	 LIS_OR2 port map( A => G442, B => G443, Z => G139 );
OR2_83:	 LIS_OR2 port map( A => G422, B => G423, Z => G532 );
OR2_84:	 LIS_OR2 port map( A => G432, B => G433, Z => G535 );
OR2_85:	 LIS_OR2 port map( A => G448, B => G449, Z => G537 );

--NAND-gates (total number: 119)
NAND2_0: LIS_NAND2 port map( A => G0, B => G2, Z => G57 );
NAND2_1: LIS_NAND2 port map( A => G1, B => G3, Z => G58 );
NAND2_2: LIS_NAND2 port map( A => G0, B => G3, Z => G76 );
NAND2_3: LIS_NAND2 port map( A => G3, B => G4, Z => G101 );
NAND2_4: LIS_NAND2 port map( A => G2, B => G4, Z => G117 );
NAND2_5: LIS_NAND2 port map( A => G1, B => G4, Z => G271 );
NAND2_6: LIS_NAND2 port map( A => G2, B => G5, Z => G97 );
NAND2_7: LIS_NAND2 port map( A => G3, B => G5, Z => G134 );
NAND2_8: LIS_NAND2 port map( A => G4, B => G6, Z => G54 );
NAND2_9: LIS_NAND2 port map( A => G6, B => G9, Z => G116 );
NAND2_10: LIS_NAND2 port map( A => G8, B => G10, Z => G71 );
NAND2_11: LIS_NAND2 port map( A => G7, B => G10, Z => G274 );
NAND2_12: LIS_NAND2 port map( A => G9, B => G11, Z => G74 );
NAND2_13: LIS_NAND2 port map( A => G8, B => G31, Z => G112 );
NAND2_14: LIS_NAND2 port map( A => G8, B => G34, Z => G245 );
NAND2_15: LIS_NAND2 port map( A => G522, B => G3, Z => G122 );
NAND2_16: LIS_NAND2 port map( A => G2, B => G524, Z => G238 );
NAND2_17: LIS_NAND2 port map( A => G527, B => G5, Z => G129 );
NAND2_18: LIS_NAND2 port map( A => G4, B => G134, Z => G240 );
NAND4_0: LIS_NAND4 port map( A => G3, B => G11, C => G35, D => G216, Z => G252 );
NAND2_19: LIS_NAND2 port map( A => G4, B => G528, Z => G77 );
NAND3_0: LIS_NAND3 port map( A => G529, B => G7, C => G30, Z => G103 );
NAND2_20: LIS_NAND2 port map( A => G527, B => G529, Z => G200 );
NAND2_21: LIS_NAND2 port map( A => G529, B => G36, Z => G248 );
NAND2_22: LIS_NAND2 port map( A => G531, B => G8, Z => G89 );
NAND2_23: LIS_NAND2 port map( A => G533, B => G10, Z => G222 );
NAND2_24: LIS_NAND2 port map( A => G7, B => G533, Z => G239 );
NAND2_25: LIS_NAND2 port map( A => G6, B => G536, Z => G235 );
NAND2_26: LIS_NAND2 port map( A => G7, B => G71, Z => G220 );
NAND2_27: LIS_NAND2 port map( A => G9, B => G538, Z => G49 );
NAND2_28: LIS_NAND2 port map( A => G543, B => G32, Z => G251 );
NAND3_1: LIS_NAND3 port map( A => G3, B => G543, C => G140, Z => G276 );
NAND2_29: LIS_NAND2 port map( A => G0, B => G99, Z => G263 );
NAND2_30: LIS_NAND2 port map( A => G527, B => G59, Z => G226 );
NAND2_31: LIS_NAND2 port map( A => G520, B => G272, Z => G210 );
NAND2_32: LIS_NAND2 port map( A => G129, B => G101, Z => G66 );
NAND2_33: LIS_NAND2 port map( A => G522, B => G135, Z => G233 );
NAND3_2: LIS_NAND3 port map( A => G122, B => G238, C => G240, Z => G104 );
NAND2_34: LIS_NAND2 port map( A => G55, B => G3, Z => G86 );
NAND2_35: LIS_NAND2 port map( A => G524, B => G55, Z => G219 );
NAND2_36: LIS_NAND2 port map( A => G302, B => G528, Z => G68 );
NAND2_37: LIS_NAND2 port map( A => G536, B => G164, Z => G232 );
NAND2_38: LIS_NAND2 port map( A => G222, B => G224, Z => G136 );
NAND2_39: LIS_NAND2 port map( A => G350, B => G235, Z => G510 );
NAND2_40: LIS_NAND2 port map( A => G316, B => G72, Z => G161 );
NAND2_41: LIS_NAND2 port map( A => G381, B => G220, Z => G100 );
NAND2_42: LIS_NAND2 port map( A => G384, B => G239, Z => G85 );
NAND3_3: LIS_NAND3 port map( A => G368, B => G275, C => G34, Z => G243 );
NAND2_43: LIS_NAND2 port map( A => G75, B => G8, Z => G63 );
NAND3_4: LIS_NAND3 port map( A => G10, B => G75, C => G201, Z => G237 );
NAND2_44: LIS_NAND2 port map( A => G286, B => G538, Z => G503 );
NAND2_45: LIS_NAND2 port map( A => G374, B => G375, Z => G56 );
NAND2_46: LIS_NAND2 port map( A => G355, B => G356, Z => G83 );
NAND2_47: LIS_NAND2 port map( A => G313, B => G314, Z => G96 );
NAND2_48: LIS_NAND2 port map( A => G332, B => G333, Z => G278 );
NAND3_5: LIS_NAND3 port map( A => G309, B => G2, C => G529, Z => G255 );
NAND3_6: LIS_NAND3 port map( A => G419, B => G420, C => G233, Z => G69 );
NAND2_49: LIS_NAND2 port map( A => G310, B => G233, Z => G512 );
NAND2_50: LIS_NAND2 port map( A => G2, B => G78, Z => G181 );
NAND3_7: LIS_NAND3 port map( A => G394, B => G395, C => G81, Z => G277 );
NAND2_51: LIS_NAND2 port map( A => G305, B => G200, Z => G151 );
NAND3_8: LIS_NAND3 port map( A => G407, B => G408, C => G409, Z => G48 );
NAND2_52: LIS_NAND2 port map( A => G227, B => G241, Z => G264 );
NAND2_53: LIS_NAND2 port map( A => G68, B => G229, Z => G208 );
NAND2_54: LIS_NAND2 port map( A => G75, B => G221, Z => G168 );
NAND2_55: LIS_NAND2 port map( A => G369, B => G370, Z => G84 );
NAND3_9: LIS_NAND3 port map( A => G464, B => G103, C => G223, Z => G258 );
NAND2_56: LIS_NAND2 port map( A => G7, B => G50, Z => G166 );
NAND2_57: LIS_NAND2 port map( A => G130, B => G225, Z => G259 );
NAND2_58: LIS_NAND2 port map( A => G292, B => G293, Z => G504 );
NAND2_59: LIS_NAND2 port map( A => G50, B => G230, Z => G217 );
NAND2_60: LIS_NAND2 port map( A => G538, B => G230, Z => G257 );
NAND3_10: LIS_NAND3 port map( A => G528, B => G529, C => G191, Z => G260 );
NAND2_61: LIS_NAND2 port map( A => G524, B => G96, Z => G266 );
NAND2_62: LIS_NAND2 port map( A => G527, B => G278, Z => G262 );
NAND2_63: LIS_NAND2 port map( A => G465, B => G263, Z => G138 );
NAND2_64: LIS_NAND2 port map( A => G4, B => G69, Z => G256 );
NAND2_65: LIS_NAND2 port map( A => G334, B => G335, Z => G82 );
NAND2_66: LIS_NAND2 port map( A => G269, B => G219, Z => G109 );
NAND2_67: LIS_NAND2 port map( A => G287, B => G524, Z => G206 );
NAND2_68: LIS_NAND2 port map( A => G521, B => G87, Z => G204 );
NAND2_69: LIS_NAND2 port map( A => G264, B => G237, Z => G53 );
NAND2_70: LIS_NAND2 port map( A => G325, B => G326, Z => G273 );
NAND2_71: LIS_NAND2 port map( A => G536, B => G84, Z => G267 );
NAND2_72: LIS_NAND2 port map( A => G389, B => G390, Z => G113 );
NAND3_11: LIS_NAND3 port map( A => G258, B => G193, C => G259, Z => G143 );
NAND2_73: LIS_NAND2 port map( A => G64, B => G275, Z => G213 );
NAND2_74: LIS_NAND2 port map( A => G260, B => G237, Z => G51 );
NAND3_12: LIS_NAND3 port map( A => G320, B => G266, C => G210, Z => G102 );
NAND3_13: LIS_NAND3 port map( A => G298, B => G299, C => G219, Z => G52 );
NAND3_14: LIS_NAND3 port map( A => G421, B => G226, C => G256, Z => G80 );
NAND2_75: LIS_NAND2 port map( A => G345, B => G204, Z => G270 );
NAND3_15: LIS_NAND3 port map( A => G261, B => G181, C => G262, Z => G94 );
NAND3_16: LIS_NAND3 port map( A => G300, B => G301, C => G181, Z => G505 );
NAND3_17: LIS_NAND3 port map( A => G11, B => G273, C => G201, Z => G249 );
NAND2_76: LIS_NAND2 port map( A => G11, B => G113, Z => G268 );
NAND2_77: LIS_NAND2 port map( A => G213, B => G217, Z => G111 );
NAND3_18: LIS_NAND3 port map( A => G296, B => G297, C => G166, Z => G534 );
NAND2_78: LIS_NAND2 port map( A => G87, B => G218, Z => G253 );
NAND3_19: LIS_NAND3 port map( A => G454, B => G455, C => G0, Z => G148 );
NAND2_79: LIS_NAND2 port map( A => G1, B => G152, Z => G254 );
NAND2_80: LIS_NAND2 port map( A => G391, B => G268, Z => G127 );
NAND3_20: LIS_NAND3 port map( A => G135, B => G55, C => G212, Z => G215 );
NAND2_81: LIS_NAND2 port map( A => G534, B => G32, Z => G62 );
NAND3_21: LIS_NAND3 port map( A => G254, B => G255, C => G208, Z => G523 );
NAND2_82: LIS_NAND2 port map( A => G318, B => G319, Z => G508 );
NAND3_22: LIS_NAND3 port map( A => G215, B => G252, C => G253, Z => G144 );
NAND2_83: LIS_NAND2 port map( A => G13, B => G523, Z => G250 );
NAND2_84: LIS_NAND2 port map( A => G523, B => G534, Z => G281 );
NAND2_85: LIS_NAND2 port map( A => G553, B => G187, Z => G171 );
NAND3_23: LIS_NAND3 port map( A => G1, B => G2, C => G141, Z => G526 );
NAND2_86: LIS_NAND2 port map( A => G46, B => G247, Z => G280 );
NAND2_87: LIS_NAND2 port map( A => G544, B => G186, Z => G246 );
NAND2_88: LIS_NAND2 port map( A => G284, B => G285, Z => G119 );
NAND2_89: LIS_NAND2 port map( A => G294, B => G295, Z => G120 );
NAND2_90: LIS_NAND2 port map( A => G525, B => G184, Z => G185 );
NAND2_91: LIS_NAND2 port map( A => G6, B => G155, Z => G159 );
NAND3_24: LIS_NAND3 port map( A => G450, B => G185, C => G246, Z => G518 );
NAND3_25: LIS_NAND3 port map( A => G243, B => G244, C => G279, Z => G542 );

--NOR-gates (total number: 50)
NOR2_0:	 LIS_NOR2 port map( A => G0, B => G4, Z => G163 );
NOR2_1:	 LIS_NOR2 port map( A => G4, B => G5, Z => G216 );
NOR2_2:	 LIS_NOR2 port map( A => G5, B => G7, Z => G169 );
NOR2_3:	 LIS_NOR2 port map( A => G7, B => G8, Z => G225 );
NOR2_4:	 LIS_NOR2 port map( A => G7, B => G11, Z => G190 );
NOR2_5:	 LIS_NOR2 port map( A => G10, B => G11, Z => G241 );
NOR2_6:	 LIS_NOR2 port map( A => G520, B => G3, Z => G198 );
NOR2_7:	 LIS_NOR2 port map( A => G521, B => G4, Z => G178 );
NOR2_8:	 LIS_NOR2 port map( A => G1, B => G522, Z => G229 );
NOR2_9:	 LIS_NOR2 port map( A => G1, B => G524, Z => G209 );
NOR2_10:	 LIS_NOR2 port map( A => G521, B => G134, Z => G195 );
NOR2_11:	 LIS_NOR2 port map( A => G522, B => G54, Z => G189 );
NOR2_12:	 LIS_NOR2 port map( A => G528, B => G54, Z => G201 );
NOR2_13:	 LIS_NOR2 port map( A => G531, B => G10, Z => G164 );
NOR2_14:	 LIS_NOR2 port map( A => G6, B => G274, Z => G211 );
NOR2_15:	 LIS_NOR2 port map( A => G12, B => G543, Z => G156 );
NOR2_16:	 LIS_NOR2 port map( A => G529, B => G122, Z => G205 );
NOR2_17:	 LIS_NOR2 port map( A => G5, B => G200, Z => G227 );
NOR2_18:	 LIS_NOR2 port map( A => G8, B => G490, Z => G230 );
NOR2_19:	 LIS_NOR2 port map( A => G9, B => G482, Z => G191 );
NOR3_0:	 LIS_NOR3 port map( A => G5, B => G540, C => G86, Z => G196 );
NOR2_20:	 LIS_NOR2 port map( A => G540, B => G232, Z => G197 );
NOR2_21:	 LIS_NOR2 port map( A => G10, B => G63, Z => G202 );
NOR2_22:	 LIS_NOR2 port map( A => G436, B => G437, Z => G502 );
NOR2_23:	 LIS_NOR2 port map( A => G528, B => G217, Z => G218 );
NOR3_1:	 LIS_NOR3 port map( A => G410, B => G411, C => G412, Z => G516 );
NOR2_24:	 LIS_NOR2 port map( A => G387, B => G388, Z => G515 );
NOR2_25:	 LIS_NOR2 port map( A => G331, B => G5, Z => G509 );
NOR2_26:	 LIS_NOR2 port map( A => G360, B => G361, Z => G513 );
NOR2_27:	 LIS_NOR2 port map( A => G330, B => G3, Z => G183 );
NOR2_28:	 LIS_NOR2 port map( A => G428, B => G429, Z => G517 );
NOR2_29:	 LIS_NOR2 port map( A => G12, B => G62, Z => G182 );
NOR4_0:	 LIS_NOR4 port map( A => G460, B => G461, C => G462, D => G463, Z => G519 );
NOR2_30:	 LIS_NOR2 port map( A => G4, B => G494, Z => G176 );
NOR2_31:	 LIS_NOR2 port map( A => G86, B => G500, Z => G175 );
NOR2_32:	 LIS_NOR2 port map( A => G13, B => G492, Z => G187 );
NOR2_33:	 LIS_NOR2 port map( A => G521, B => G281, Z => G158 );
NOR2_34:	 LIS_NOR2 port map( A => G281, B => G271, Z => G194 );
NOR2_35:	 LIS_NOR2 port map( A => G13, B => G483, Z => G157 );
NOR3_2:	 LIS_NOR3 port map( A => G315, B => G12, C => G487, Z => G507 );
NOR2_36:	 LIS_NOR2 port map( A => G282, B => G501, Z => G186 );
NOR4_1:	 LIS_NOR4 port map( A => G471, B => G472, C => G473, D => G474, Z => G247 );
NOR2_37:	 LIS_NOR2 port map( A => G541, B => G280, Z => G179 );
NOR2_38:	 LIS_NOR2 port map( A => G543, B => G493, Z => G188 );
NOR2_39:	 LIS_NOR2 port map( A => G12, B => G488, Z => G154 );
NOR3_3:	 LIS_NOR3 port map( A => G541, B => G13, C => G499, Z => G184 );
NOR2_40:	 LIS_NOR2 port map( A => G311, B => G312, Z => G506 );
NOR2_41:	 LIS_NOR2 port map( A => G13, B => G480, Z => G155 );
NOR2_42:	 LIS_NOR2 port map( A => G185, B => G498, Z => G162 );
NOR3_4:	 LIS_NOR3 port map( A => G372, B => G373, C => G478, Z => G514 );

end architecture;
